module bgf_rom
	(
		input wire clk,
		input wire [7:0] row,
		input wire [7:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [7:0] row_reg;
	reg [7:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin
		if(({row_reg, col_reg}>=16'b0000000000000000) && ({row_reg, col_reg}<16'b0000000000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000000001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000000001101) && ({row_reg, col_reg}<16'b0000000000001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000000000001111) && ({row_reg, col_reg}<16'b0000000000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000000010001) && ({row_reg, col_reg}<16'b0000000000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000000000100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000000100110) && ({row_reg, col_reg}<16'b0000000000101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000000101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000000101010) && ({row_reg, col_reg}<16'b0000000000101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000000101101) && ({row_reg, col_reg}<16'b0000000000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000000110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000000110010) && ({row_reg, col_reg}<16'b0000000000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000000110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000000000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000000000110111) && ({row_reg, col_reg}<16'b0000000000111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000000000111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000000000111010) && ({row_reg, col_reg}<16'b0000000000111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000000111100) && ({row_reg, col_reg}<16'b0000000000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000000000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000000111111) && ({row_reg, col_reg}<16'b0000000001000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000001000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000000001000100) && ({row_reg, col_reg}<16'b0000000001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000001000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000000001000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000001001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000001001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000000001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000001001011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0000000001001100) && ({row_reg, col_reg}<16'b0000000001001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000000001001110) && ({row_reg, col_reg}<16'b0000000001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000001010100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0000000001010101) && ({row_reg, col_reg}<16'b0000000001010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000000001010111) && ({row_reg, col_reg}<16'b0000000001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000001011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000000001100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000001100001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000000001100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000000001100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000001100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000000001100101) && ({row_reg, col_reg}<16'b0000000001100111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000000001100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000001101000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000000001101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000000001101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0000000001101011) && ({row_reg, col_reg}<16'b0000000001101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000000001101101) && ({row_reg, col_reg}<16'b0000000001101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000001101111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000000001110000)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0000000001110001) && ({row_reg, col_reg}<16'b0000000001110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000001110011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000000001110100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000000001110101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000000001110110) && ({row_reg, col_reg}<16'b0000000001111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000001111000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000000001111001) && ({row_reg, col_reg}<16'b0000000001111100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0000000001111100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0000000001111101) && ({row_reg, col_reg}<16'b0000000001111111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0000000001111111)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0000000010000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000000010000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000010000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000000010000011) && ({row_reg, col_reg}<16'b0000000010000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000010000101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000010000110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000000010000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000000010001000) && ({row_reg, col_reg}<16'b0000000010001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000010001100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000000010001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000010001110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000000010001111) && ({row_reg, col_reg}<16'b0000000010010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000010010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000000010010011) && ({row_reg, col_reg}<16'b0000000010010101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000000010010101) && ({row_reg, col_reg}<16'b0000000010010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000000010010111) && ({row_reg, col_reg}<16'b0000000010011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000010011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000000010011101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000000010011110) && ({row_reg, col_reg}<16'b0000000010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000010100011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0000000010100100) && ({row_reg, col_reg}<16'b0000000010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000000010100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0000000010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000000010101000) && ({row_reg, col_reg}<16'b0000000010101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000000010101011) && ({row_reg, col_reg}<16'b0000000010110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000000010110001) && ({row_reg, col_reg}<16'b0000000010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000000010110011) && ({row_reg, col_reg}<16'b0000000010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000000010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000000010111001) && ({row_reg, col_reg}<16'b0000000010111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000010111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000000010111111) && ({row_reg, col_reg}<16'b0000000011000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000011000010) && ({row_reg, col_reg}<16'b0000000011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000000011000100) && ({row_reg, col_reg}<16'b0000000011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000011000110) && ({row_reg, col_reg}<16'b0000000011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000011001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000000011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000000011001100) && ({row_reg, col_reg}<16'b0000000011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000000011001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000000011001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000011010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000011010001) && ({row_reg, col_reg}<16'b0000000011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000000011110000) && ({row_reg, col_reg}<16'b0000000011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000000011110011) && ({row_reg, col_reg}<16'b0000000011110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000011110110) && ({row_reg, col_reg}<16'b0000000011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000000011111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000000011111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000011111011) && ({row_reg, col_reg}<16'b0000000011111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0000000011111110) && ({row_reg, col_reg}<16'b0000000100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000100000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000000100000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000000100000011) && ({row_reg, col_reg}<16'b0000000100001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000100001011) && ({row_reg, col_reg}<16'b0000000100001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000000100001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000000100001110) && ({row_reg, col_reg}<16'b0000000100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000100010010) && ({row_reg, col_reg}<16'b0000000100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000000100100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000100100110) && ({row_reg, col_reg}<16'b0000000100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000100101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000100101010) && ({row_reg, col_reg}<16'b0000000100101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000100101101) && ({row_reg, col_reg}<16'b0000000100110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000100110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000100110010) && ({row_reg, col_reg}<16'b0000000100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000100110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000000100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000100110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000000100110111) && ({row_reg, col_reg}<16'b0000000100111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000000100111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000100111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000100111011) && ({row_reg, col_reg}<16'b0000000100111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000000100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000100111111) && ({row_reg, col_reg}<16'b0000000101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000101000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000000101000100) && ({row_reg, col_reg}<16'b0000000101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000000101000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000101001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000000101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000000101001100) && ({row_reg, col_reg}<16'b0000000101001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000000101001110) && ({row_reg, col_reg}<16'b0000000101010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000101010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000000101010110) && ({row_reg, col_reg}<16'b0000000101011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000101011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000000101100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000101100001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000000101100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000000101100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000000101100100) && ({row_reg, col_reg}<16'b0000000101101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000101101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000000101101001) && ({row_reg, col_reg}<16'b0000000101101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000000101101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000000101101100) && ({row_reg, col_reg}<16'b0000000101101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000000101101110) && ({row_reg, col_reg}<16'b0000000101110001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000000101110001) && ({row_reg, col_reg}<16'b0000000101110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000101110011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000000101110100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000000101110101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000000101110110) && ({row_reg, col_reg}<16'b0000000101111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000000101111000) && ({row_reg, col_reg}<16'b0000000101111010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000000101111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000101111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000101111100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0000000101111101) && ({row_reg, col_reg}<16'b0000000101111111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0000000101111111) && ({row_reg, col_reg}<16'b0000000110000001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000000110000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000110000010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000000110000011) && ({row_reg, col_reg}<16'b0000000110000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000110000101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000110000110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000000110000111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000000110001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000000110001001) && ({row_reg, col_reg}<16'b0000000110001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000110001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000110001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000110001110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000000110001111) && ({row_reg, col_reg}<16'b0000000110010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000000110010010) && ({row_reg, col_reg}<16'b0000000110010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000110010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000000110010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000110011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000000110011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000110011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000000110011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000000110011110) && ({row_reg, col_reg}<16'b0000000110100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000000110100011) && ({row_reg, col_reg}<16'b0000000110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000000110100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0000000110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000000110101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000000110101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000000110101011) && ({row_reg, col_reg}<16'b0000000110110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000110110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000000110110001) && ({row_reg, col_reg}<16'b0000000110110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000000110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000000110110100) && ({row_reg, col_reg}<16'b0000000110110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000000110110110) && ({row_reg, col_reg}<16'b0000000110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000000110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000000110111001) && ({row_reg, col_reg}<16'b0000000110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000000110111101) && ({row_reg, col_reg}<16'b0000000110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000000110111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000111000010) && ({row_reg, col_reg}<16'b0000000111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000000111000100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000111000101) && ({row_reg, col_reg}<16'b0000000111001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000111001010) && ({row_reg, col_reg}<16'b0000000111001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000111001100) && ({row_reg, col_reg}<16'b0000000111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000111001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000111001111) && ({row_reg, col_reg}<16'b0000000111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000111010001) && ({row_reg, col_reg}<16'b0000000111110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000000111110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000111110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000000111110010) && ({row_reg, col_reg}<16'b0000000111110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000111110110) && ({row_reg, col_reg}<16'b0000000111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000000111111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000000111111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000111111011) && ({row_reg, col_reg}<16'b0000000111111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0000000111111110) && ({row_reg, col_reg}<16'b0000001000000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000001000000001)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==16'b0000001000000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000001000000011) && ({row_reg, col_reg}<16'b0000001000000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001000000101) && ({row_reg, col_reg}<16'b0000001000001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001000001011) && ({row_reg, col_reg}<16'b0000001000001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000001000001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000001000001110) && ({row_reg, col_reg}<16'b0000001000010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000001000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001000010010) && ({row_reg, col_reg}<16'b0000001000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000001000100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001000100110) && ({row_reg, col_reg}<16'b0000001000101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000001000101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001000101010) && ({row_reg, col_reg}<16'b0000001000101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001000101101) && ({row_reg, col_reg}<16'b0000001000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001000110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001000110010) && ({row_reg, col_reg}<16'b0000001000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001000110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000001000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000001000110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001000111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000001000111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000001000111010) && ({row_reg, col_reg}<16'b0000001000111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001000111100) && ({row_reg, col_reg}<16'b0000001000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000001000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001000111111) && ({row_reg, col_reg}<16'b0000001001000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000001001000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000001001000100) && ({row_reg, col_reg}<16'b0000001001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001001000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000001001000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001001001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000001001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000001001001100) && ({row_reg, col_reg}<16'b0000001001001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000001001001110) && ({row_reg, col_reg}<16'b0000001001010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001001010101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000001001010110) && ({row_reg, col_reg}<16'b0000001001011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001001011010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000001001011011) && ({row_reg, col_reg}<16'b0000001001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001001011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000001001100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001001100001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000001001100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000001001100011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0000001001100100) && ({row_reg, col_reg}<16'b0000001001101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001001101001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000001001101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000001001101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000001001101100) && ({row_reg, col_reg}<16'b0000001001101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000001001101110) && ({row_reg, col_reg}<16'b0000001001110001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000001001110001) && ({row_reg, col_reg}<16'b0000001001110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001001110011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000001001110100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001001110101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000001001110110) && ({row_reg, col_reg}<16'b0000001001111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001001111000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000001001111001) && ({row_reg, col_reg}<16'b0000001001111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000001001111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001001111100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0000001001111101) && ({row_reg, col_reg}<16'b0000001010000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0000001010000000) && ({row_reg, col_reg}<16'b0000001010000010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001010000010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000001010000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001010000100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000001010000101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001010000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001010000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001010001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000001010001001) && ({row_reg, col_reg}<16'b0000001010001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001010001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001010001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001010001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001010010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000001010010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000001010010010) && ({row_reg, col_reg}<16'b0000001010010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001010010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000001010010111) && ({row_reg, col_reg}<16'b0000001010011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001010011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001010011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000001010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000001010011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000001010011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000001010011111) && ({row_reg, col_reg}<16'b0000001010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000001010100011) && ({row_reg, col_reg}<16'b0000001010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000001010100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0000001010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000001010101000) && ({row_reg, col_reg}<16'b0000001010101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000001010101011) && ({row_reg, col_reg}<16'b0000001010101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001010101101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000001010101110) && ({row_reg, col_reg}<16'b0000001010110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000001010110001) && ({row_reg, col_reg}<16'b0000001010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000001010110100) && ({row_reg, col_reg}<16'b0000001010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000001010110110) && ({row_reg, col_reg}<16'b0000001010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000001010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000001010111001) && ({row_reg, col_reg}<16'b0000001010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000001010111100)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==16'b0000001010111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000001010111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000001010111111) && ({row_reg, col_reg}<16'b0000001011000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001011000010) && ({row_reg, col_reg}<16'b0000001011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000001011000100) && ({row_reg, col_reg}<16'b0000001011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001011000110) && ({row_reg, col_reg}<16'b0000001011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001011001010) && ({row_reg, col_reg}<16'b0000001011001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001011001100) && ({row_reg, col_reg}<16'b0000001011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001011001111) && ({row_reg, col_reg}<16'b0000001011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001011010001) && ({row_reg, col_reg}<16'b0000001011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000001011110000) && ({row_reg, col_reg}<16'b0000001011110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000001011110010) && ({row_reg, col_reg}<16'b0000001011110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001011110110) && ({row_reg, col_reg}<16'b0000001011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000001011111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000001011111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001011111011) && ({row_reg, col_reg}<16'b0000001011111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0000001011111110) && ({row_reg, col_reg}<16'b0000001100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000001100000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000001100000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000001100000100) && ({row_reg, col_reg}<16'b0000001100000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001100000110) && ({row_reg, col_reg}<16'b0000001100001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001100001011) && ({row_reg, col_reg}<16'b0000001100001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001100001101) && ({row_reg, col_reg}<16'b0000001100001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000001100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000001100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001100010010) && ({row_reg, col_reg}<16'b0000001100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000001100100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001100100110) && ({row_reg, col_reg}<16'b0000001100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000001100101000) && ({row_reg, col_reg}<16'b0000001100101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001100101010) && ({row_reg, col_reg}<16'b0000001100101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000001100101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000001100101110) && ({row_reg, col_reg}<16'b0000001100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001100110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000001100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000001100110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000001100111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000001100111001) && ({row_reg, col_reg}<16'b0000001100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000001100111011) && ({row_reg, col_reg}<16'b0000001100111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001100111111) && ({row_reg, col_reg}<16'b0000001101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000001101000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000001101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001101000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000001101000111) && ({row_reg, col_reg}<16'b0000001101001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000001101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000001101001010) && ({row_reg, col_reg}<16'b0000001101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000001101001100) && ({row_reg, col_reg}<16'b0000001101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000001101001111) && ({row_reg, col_reg}<16'b0000001101011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001101011011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000001101011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001101011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001101011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000001101100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001101100001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000001101100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000001101100011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000001101100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000001101100101) && ({row_reg, col_reg}<16'b0000001101100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000001101100111) && ({row_reg, col_reg}<16'b0000001101101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000001101101001) && ({row_reg, col_reg}<16'b0000001101101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000001101101011) && ({row_reg, col_reg}<16'b0000001101110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000001101110000)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0000001101110001) && ({row_reg, col_reg}<16'b0000001101110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000001101110011) && ({row_reg, col_reg}<16'b0000001101110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000001101110101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000001101110110) && ({row_reg, col_reg}<16'b0000001101111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001101111000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000001101111001) && ({row_reg, col_reg}<16'b0000001101111100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000001101111100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000001101111101) && ({row_reg, col_reg}<16'b0000001101111111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001101111111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0000001110000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0000001110000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001110000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000001110000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000001110000100) && ({row_reg, col_reg}<16'b0000001110000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001110000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000001110000111) && ({row_reg, col_reg}<16'b0000001110001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001110001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001110001101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000001110001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001110001111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000001110010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000001110010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000001110010010) && ({row_reg, col_reg}<16'b0000001110010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001110010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000001110010111) && ({row_reg, col_reg}<16'b0000001110011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001110011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000001110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000001110011101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0000001110011110) && ({row_reg, col_reg}<16'b0000001110100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000001110100000) && ({row_reg, col_reg}<16'b0000001110100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000001110100011) && ({row_reg, col_reg}<16'b0000001110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000001110100110) && ({row_reg, col_reg}<16'b0000001110101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000001110101001) && ({row_reg, col_reg}<16'b0000001110101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001110101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000001110101100) && ({row_reg, col_reg}<16'b0000001110101110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000001110101110) && ({row_reg, col_reg}<16'b0000001110110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000001110110001) && ({row_reg, col_reg}<16'b0000001110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000001110110100) && ({row_reg, col_reg}<16'b0000001110110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000001110110110) && ({row_reg, col_reg}<16'b0000001110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000001110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000001110111001) && ({row_reg, col_reg}<16'b0000001110111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000001110111100)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==16'b0000001110111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000001110111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000001110111111) && ({row_reg, col_reg}<16'b0000001111000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000001111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001111000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000001111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000001111000100) && ({row_reg, col_reg}<16'b0000001111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001111000110) && ({row_reg, col_reg}<16'b0000001111001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001111001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000001111001100) && ({row_reg, col_reg}<16'b0000001111001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001111001111) && ({row_reg, col_reg}<16'b0000001111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001111010001) && ({row_reg, col_reg}<16'b0000001111110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000001111110000) && ({row_reg, col_reg}<16'b0000001111110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000001111110010) && ({row_reg, col_reg}<16'b0000001111111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000001111111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001111111011) && ({row_reg, col_reg}<16'b0000001111111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000001111111110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0000001111111111) && ({row_reg, col_reg}<16'b0000010000000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010000000011) && ({row_reg, col_reg}<16'b0000010000000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010000000111) && ({row_reg, col_reg}<16'b0000010000001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010000001011) && ({row_reg, col_reg}<16'b0000010000001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010000001101) && ({row_reg, col_reg}<16'b0000010000001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000010000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010000010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000010000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010000010010) && ({row_reg, col_reg}<16'b0000010000100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000010000100100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010000100101) && ({row_reg, col_reg}<16'b0000010000100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010000100111) && ({row_reg, col_reg}<16'b0000010000101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000010000101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010000101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010000101011) && ({row_reg, col_reg}<16'b0000010000101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000010000101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000010000101110) && ({row_reg, col_reg}<16'b0000010000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010000110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000010000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000010000110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000010000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010000111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000010000111010) && ({row_reg, col_reg}<16'b0000010000111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010000111111) && ({row_reg, col_reg}<16'b0000010001000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000010001000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000010001000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010001000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000010001001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000010001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000010001001010) && ({row_reg, col_reg}<16'b0000010001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010001001100) && ({row_reg, col_reg}<16'b0000010001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000010001001111) && ({row_reg, col_reg}<16'b0000010001010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010001010111) && ({row_reg, col_reg}<16'b0000010001011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000010001011010) && ({row_reg, col_reg}<16'b0000010001011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010001011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010001011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010001011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000010001100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010001100001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000010001100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000010001100011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000010001100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000010001100101) && ({row_reg, col_reg}<16'b0000010001100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000010001100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010001101000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000010001101001) && ({row_reg, col_reg}<16'b0000010001101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010001101011) && ({row_reg, col_reg}<16'b0000010001110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000010001110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000010001110001) && ({row_reg, col_reg}<16'b0000010001110100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000010001110100) && ({row_reg, col_reg}<16'b0000010001110110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000010001110110) && ({row_reg, col_reg}<16'b0000010001111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010001111000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000010001111001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000010001111010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000010001111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000010001111100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000010001111101) && ({row_reg, col_reg}<16'b0000010010000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010010000000)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0000010010000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010010000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000010010000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000010010000100) && ({row_reg, col_reg}<16'b0000010010000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010010000110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000010010000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000010010001000) && ({row_reg, col_reg}<16'b0000010010001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010010001100) && ({row_reg, col_reg}<16'b0000010010001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010010001111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000010010010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010010010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000010010010010) && ({row_reg, col_reg}<16'b0000010010010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010010010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000010010010110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0000010010010111) && ({row_reg, col_reg}<16'b0000010010011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010010011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000010010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000010010011101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000010010011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010010011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010010100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000010010100001) && ({row_reg, col_reg}<16'b0000010010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010010100011) && ({row_reg, col_reg}<16'b0000010010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000010010100110) && ({row_reg, col_reg}<16'b0000010010101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000010010101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000010010101010) && ({row_reg, col_reg}<16'b0000010010101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010010101100) && ({row_reg, col_reg}<16'b0000010010110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000010010110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010010110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010010110010)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}==16'b0000010010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000010010110100) && ({row_reg, col_reg}<16'b0000010010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000010010110110) && ({row_reg, col_reg}<16'b0000010010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000010010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010010111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000010010111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010010111011) && ({row_reg, col_reg}<16'b0000010010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000010010111101) && ({row_reg, col_reg}<16'b0000010010111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000010010111111) && ({row_reg, col_reg}<16'b0000010011000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000010011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010011000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000010011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000010011000100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000010011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000010011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010011000111) && ({row_reg, col_reg}<16'b0000010011001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010011001011) && ({row_reg, col_reg}<16'b0000010011001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010011001101) && ({row_reg, col_reg}<16'b0000010011001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000010011001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000010011010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010011010001) && ({row_reg, col_reg}<16'b0000010011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000010011110000) && ({row_reg, col_reg}<16'b0000010011110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000010011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000010011110011) && ({row_reg, col_reg}<16'b0000010011110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000010011110110)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=16'b0000010011110111) && ({row_reg, col_reg}<16'b0000010011111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000010011111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010011111011) && ({row_reg, col_reg}<16'b0000010011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000010011111110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0000010011111111) && ({row_reg, col_reg}<16'b0000010100000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000010100000011) && ({row_reg, col_reg}<16'b0000010100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010100000101) && ({row_reg, col_reg}<16'b0000010100001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010100001000) && ({row_reg, col_reg}<16'b0000010100001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010100001011) && ({row_reg, col_reg}<16'b0000010100001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010100001101) && ({row_reg, col_reg}<16'b0000010100001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000010100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010100010000) && ({row_reg, col_reg}<16'b0000010100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000010100010010) && ({row_reg, col_reg}<16'b0000010100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000010100100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000010100100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010100100111) && ({row_reg, col_reg}<16'b0000010100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000010100101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010100101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010100101011) && ({row_reg, col_reg}<16'b0000010100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000010100101101) && ({row_reg, col_reg}<16'b0000010100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010100110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000010100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010100110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000010100110111) && ({row_reg, col_reg}<16'b0000010100111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010100111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000010100111010) && ({row_reg, col_reg}<16'b0000010100111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010100111100) && ({row_reg, col_reg}<16'b0000010100111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000010100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010100111111) && ({row_reg, col_reg}<16'b0000010101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000010101000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000010101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000010101000111) && ({row_reg, col_reg}<16'b0000010101001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000010101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010101001011) && ({row_reg, col_reg}<16'b0000010101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010101001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010101010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000010101010001) && ({row_reg, col_reg}<16'b0000010101010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010101010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010101011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000010101011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000010101011010) && ({row_reg, col_reg}<16'b0000010101011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010101011111) && ({row_reg, col_reg}<16'b0000010101100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010101100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010101100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000010101100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010101100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010101100101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000010101100110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000010101100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000010101101000) && ({row_reg, col_reg}<16'b0000010101101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000010101101011) && ({row_reg, col_reg}<16'b0000010101101111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000010101101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010101110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000010101110001) && ({row_reg, col_reg}<16'b0000010101110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010101110101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000010101110110) && ({row_reg, col_reg}<16'b0000010101111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010101111000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000010101111001) && ({row_reg, col_reg}<16'b0000010101111100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000010101111100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000010101111101) && ({row_reg, col_reg}<16'b0000010110000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010110000000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000010110000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010110000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000010110000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010110000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010110000101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000010110000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010110000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010110001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010110001001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000010110001010) && ({row_reg, col_reg}<16'b0000010110001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010110001100) && ({row_reg, col_reg}<16'b0000010110001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010110001111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000010110010000) && ({row_reg, col_reg}<16'b0000010110010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010110010010) && ({row_reg, col_reg}<16'b0000010110010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010110010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000010110010110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0000010110010111) && ({row_reg, col_reg}<16'b0000010110011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010110011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000010110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000010110011101) && ({row_reg, col_reg}<16'b0000010110100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010110100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000010110100001) && ({row_reg, col_reg}<16'b0000010110100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010110100011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0000010110100100) && ({row_reg, col_reg}<16'b0000010110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000010110100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0000010110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010110101000) && ({row_reg, col_reg}<16'b0000010110101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010110101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010110101011) && ({row_reg, col_reg}<16'b0000010110110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000010110110000) && ({row_reg, col_reg}<16'b0000010110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010110110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000010110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000010110110110) && ({row_reg, col_reg}<16'b0000010110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000010110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010110111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000010110111010) && ({row_reg, col_reg}<16'b0000010110111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000010110111110) && ({row_reg, col_reg}<16'b0000010111000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000010111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010111000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000010111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000010111000100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000010111000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000010111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010111000111) && ({row_reg, col_reg}<16'b0000010111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010111001001) && ({row_reg, col_reg}<16'b0000010111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000010111001011) && ({row_reg, col_reg}<16'b0000010111001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010111001101) && ({row_reg, col_reg}<16'b0000010111001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000010111001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000010111010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010111010001) && ({row_reg, col_reg}<16'b0000010111110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000010111110000) && ({row_reg, col_reg}<16'b0000010111110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000010111110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010111110011) && ({row_reg, col_reg}<16'b0000010111110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010111110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010111110110) && ({row_reg, col_reg}<16'b0000010111111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000010111111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010111111011) && ({row_reg, col_reg}<16'b0000010111111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000010111111110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}==16'b0000010111111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011000000000) && ({row_reg, col_reg}<16'b0000011000000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000011000000100) && ({row_reg, col_reg}<16'b0000011000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011000000110) && ({row_reg, col_reg}<16'b0000011000001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011000001001) && ({row_reg, col_reg}<16'b0000011000001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011000001011) && ({row_reg, col_reg}<16'b0000011000001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011000001101) && ({row_reg, col_reg}<16'b0000011000001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000011000001111) && ({row_reg, col_reg}<16'b0000011000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011000010010) && ({row_reg, col_reg}<16'b0000011000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000011000100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000011000100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011000100111) && ({row_reg, col_reg}<16'b0000011000101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000011000101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011000101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011000101011) && ({row_reg, col_reg}<16'b0000011000101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000011000101101) && ({row_reg, col_reg}<16'b0000011000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011000110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000011000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000011000110111) && ({row_reg, col_reg}<16'b0000011000111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000011000111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000011000111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011000111011) && ({row_reg, col_reg}<16'b0000011000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000011000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011000111111) && ({row_reg, col_reg}<16'b0000011001000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000011001000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000011001000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000011001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011001000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000011001000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011001001000) && ({row_reg, col_reg}<16'b0000011001001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000011001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000011001001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000011001001101) && ({row_reg, col_reg}<16'b0000011001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000011001001111) && ({row_reg, col_reg}<16'b0000011001010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000011001010111) && ({row_reg, col_reg}<16'b0000011001011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000011001011010) && ({row_reg, col_reg}<16'b0000011001011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011001011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000011001011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000011001011111) && ({row_reg, col_reg}<16'b0000011001100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011001100001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000011001100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000011001100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011001100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000011001100101) && ({row_reg, col_reg}<16'b0000011001100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011001100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000011001101000) && ({row_reg, col_reg}<16'b0000011001101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000011001101011) && ({row_reg, col_reg}<16'b0000011001101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000011001101101) && ({row_reg, col_reg}<16'b0000011001101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011001101111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000011001110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000011001110001) && ({row_reg, col_reg}<16'b0000011001111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011001111000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000011001111001) && ({row_reg, col_reg}<16'b0000011001111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000011001111100) && ({row_reg, col_reg}<16'b0000011001111110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000011001111110) && ({row_reg, col_reg}<16'b0000011010000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011010000000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000011010000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011010000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011010000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000011010000100) && ({row_reg, col_reg}<16'b0000011010000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011010000110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000011010000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011010001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011010001001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000011010001010) && ({row_reg, col_reg}<16'b0000011010001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000011010001100) && ({row_reg, col_reg}<16'b0000011010001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011010001111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000011010010000) && ({row_reg, col_reg}<16'b0000011010010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000011010010010) && ({row_reg, col_reg}<16'b0000011010010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011010010100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000011010010101) && ({row_reg, col_reg}<16'b0000011010010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000011010010111) && ({row_reg, col_reg}<16'b0000011010011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011010011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000011010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000011010011101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000011010011110) && ({row_reg, col_reg}<16'b0000011010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000011010100011) && ({row_reg, col_reg}<16'b0000011010100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000011010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000011010101001) && ({row_reg, col_reg}<16'b0000011010101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000011010101011) && ({row_reg, col_reg}<16'b0000011010110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000011010110000) && ({row_reg, col_reg}<16'b0000011010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000011010110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000011010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011010110110) && ({row_reg, col_reg}<16'b0000011010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000011010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000011010111001) && ({row_reg, col_reg}<16'b0000011010111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000011010111011) && ({row_reg, col_reg}<16'b0000011010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011010111101) && ({row_reg, col_reg}<16'b0000011010111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011010111111) && ({row_reg, col_reg}<16'b0000011011000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000011011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011011000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000011011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000011011000100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000011011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000011011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011011000111) && ({row_reg, col_reg}<16'b0000011011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011011001001) && ({row_reg, col_reg}<16'b0000011011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011011001011) && ({row_reg, col_reg}<16'b0000011011001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011011001101) && ({row_reg, col_reg}<16'b0000011011001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000011011001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011011010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011011010001) && ({row_reg, col_reg}<16'b0000011011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000011011110000) && ({row_reg, col_reg}<16'b0000011011110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011011110010) && ({row_reg, col_reg}<16'b0000011011110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011011110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000011011110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011011110111) && ({row_reg, col_reg}<16'b0000011011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011011111001) && ({row_reg, col_reg}<16'b0000011011111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011011111011) && ({row_reg, col_reg}<16'b0000011011111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0000011011111110) && ({row_reg, col_reg}<16'b0000011100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011100000000) && ({row_reg, col_reg}<16'b0000011100000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000011100000101) && ({row_reg, col_reg}<16'b0000011100000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011100000111) && ({row_reg, col_reg}<16'b0000011100001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011100001010) && ({row_reg, col_reg}<16'b0000011100001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011100001100) && ({row_reg, col_reg}<16'b0000011100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011100001111) && ({row_reg, col_reg}<16'b0000011100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011100010010) && ({row_reg, col_reg}<16'b0000011100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000011100100110) && ({row_reg, col_reg}<16'b0000011100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011100101001) && ({row_reg, col_reg}<16'b0000011100101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000011100101101) && ({row_reg, col_reg}<16'b0000011100110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011100110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011100110010) && ({row_reg, col_reg}<16'b0000011100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011100110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000011100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000011100110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011100111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000011100111001) && ({row_reg, col_reg}<16'b0000011100111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000011100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011100111111) && ({row_reg, col_reg}<16'b0000011101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000011101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000011101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000011101000111) && ({row_reg, col_reg}<16'b0000011101001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011101001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000011101001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000011101001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000011101001100) && ({row_reg, col_reg}<16'b0000011101001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000011101001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000011101001111) && ({row_reg, col_reg}<16'b0000011101010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000011101010111) && ({row_reg, col_reg}<16'b0000011101011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000011101011010) && ({row_reg, col_reg}<16'b0000011101011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000011101011111) && ({row_reg, col_reg}<16'b0000011101100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011101100001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000011101100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000011101100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011101100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000011101100101) && ({row_reg, col_reg}<16'b0000011101100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011101100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000011101101000) && ({row_reg, col_reg}<16'b0000011101101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000011101101011) && ({row_reg, col_reg}<16'b0000011101101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000011101101101) && ({row_reg, col_reg}<16'b0000011101110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000011101110001) && ({row_reg, col_reg}<16'b0000011101111001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011101111001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000011101111010) && ({row_reg, col_reg}<16'b0000011101111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011101111101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0000011101111110) && ({row_reg, col_reg}<16'b0000011110000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011110000000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000011110000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011110000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011110000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000011110000100) && ({row_reg, col_reg}<16'b0000011110000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011110000110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000011110000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011110001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011110001001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000011110001010) && ({row_reg, col_reg}<16'b0000011110001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011110001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011110001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011110001110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000011110001111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000011110010000) && ({row_reg, col_reg}<16'b0000011110010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011110010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011110010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000011110010100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0000011110010101) && ({row_reg, col_reg}<16'b0000011110010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000011110010111) && ({row_reg, col_reg}<16'b0000011110011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011110011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000011110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000011110011101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000011110011110) && ({row_reg, col_reg}<16'b0000011110100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000011110100011) && ({row_reg, col_reg}<16'b0000011110100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000011110100111) && ({row_reg, col_reg}<16'b0000011110101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000011110101100) && ({row_reg, col_reg}<16'b0000011110110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000011110110000) && ({row_reg, col_reg}<16'b0000011110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000011110110100) && ({row_reg, col_reg}<16'b0000011110110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000011110110110) && ({row_reg, col_reg}<16'b0000011110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0000011110111000) && ({row_reg, col_reg}<16'b0000011110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000011110111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000011110111011) && ({row_reg, col_reg}<16'b0000011110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011110111101) && ({row_reg, col_reg}<16'b0000011110111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011110111111) && ({row_reg, col_reg}<16'b0000011111000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000011111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011111000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000011111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000011111000100) && ({row_reg, col_reg}<16'b0000011111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011111000110) && ({row_reg, col_reg}<16'b0000011111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011111001001) && ({row_reg, col_reg}<16'b0000011111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011111001011) && ({row_reg, col_reg}<16'b0000011111001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011111001110) && ({row_reg, col_reg}<16'b0000011111010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011111010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011111010001) && ({row_reg, col_reg}<16'b0000011111110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000011111110000) && ({row_reg, col_reg}<16'b0000011111110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011111110010) && ({row_reg, col_reg}<16'b0000011111110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011111110111) && ({row_reg, col_reg}<16'b0000011111111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000011111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000011111111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011111111011) && ({row_reg, col_reg}<16'b0000011111111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000011111111110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}==16'b0000011111111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100000000000) && ({row_reg, col_reg}<16'b0000100000000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000100000000110) && ({row_reg, col_reg}<16'b0000100000001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100000001000) && ({row_reg, col_reg}<16'b0000100000001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000100000001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100000001100) && ({row_reg, col_reg}<16'b0000100000010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100000010000) && ({row_reg, col_reg}<16'b0000100000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100000010010) && ({row_reg, col_reg}<16'b0000100000100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000100000100110) && ({row_reg, col_reg}<16'b0000100000101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100000101010) && ({row_reg, col_reg}<16'b0000100000101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100000101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000100000101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100000101110) && ({row_reg, col_reg}<16'b0000100000110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000100000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100000110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100000110010) && ({row_reg, col_reg}<16'b0000100000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100000110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000100000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100000110111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000100000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100000111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000100000111010) && ({row_reg, col_reg}<16'b0000100000111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100000111100) && ({row_reg, col_reg}<16'b0000100000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000100000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100000111111) && ({row_reg, col_reg}<16'b0000100001000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000100001000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100001000110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0000100001000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000100001001000) && ({row_reg, col_reg}<16'b0000100001001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000100001001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100001001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000100001001100) && ({row_reg, col_reg}<16'b0000100001001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000100001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100001001111) && ({row_reg, col_reg}<16'b0000100001010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100001010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100001011000) && ({row_reg, col_reg}<16'b0000100001011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000100001011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100001011011) && ({row_reg, col_reg}<16'b0000100001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000100001011111) && ({row_reg, col_reg}<16'b0000100001100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100001100001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000100001100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000100001100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100001100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000100001100101) && ({row_reg, col_reg}<16'b0000100001100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000100001100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100001101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100001101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100001101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0000100001101011) && ({row_reg, col_reg}<16'b0000100001101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000100001101101) && ({row_reg, col_reg}<16'b0000100001110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000100001110001) && ({row_reg, col_reg}<16'b0000100001111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100001111010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000100001111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100001111100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0000100001111101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0000100001111110) && ({row_reg, col_reg}<16'b0000100010000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100010000000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000100010000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100010000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100010000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100010000100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000100010000101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000100010000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100010000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100010001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100010001001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000100010001010) && ({row_reg, col_reg}<16'b0000100010001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000100010001101) && ({row_reg, col_reg}<16'b0000100010001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100010001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000100010010000) && ({row_reg, col_reg}<16'b0000100010010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100010010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100010010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000100010010100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0000100010010101) && ({row_reg, col_reg}<16'b0000100010010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000100010010111) && ({row_reg, col_reg}<16'b0000100010011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100010011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000100010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000100010011101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000100010011110) && ({row_reg, col_reg}<16'b0000100010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000100010100011) && ({row_reg, col_reg}<16'b0000100010100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000100010100111) && ({row_reg, col_reg}<16'b0000100010101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000100010101100) && ({row_reg, col_reg}<16'b0000100010110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000100010110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100010110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100010110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100010110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000100010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000100010110110) && ({row_reg, col_reg}<16'b0000100010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0000100010111000) && ({row_reg, col_reg}<16'b0000100010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100010111010) && ({row_reg, col_reg}<16'b0000100010111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000100010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100010111101) && ({row_reg, col_reg}<16'b0000100010111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100011000000) && ({row_reg, col_reg}<16'b0000100011000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100011000010) && ({row_reg, col_reg}<16'b0000100011000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000100011000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100011000110) && ({row_reg, col_reg}<16'b0000100011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100011001011) && ({row_reg, col_reg}<16'b0000100011001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100011001111) && ({row_reg, col_reg}<16'b0000100011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100011010001) && ({row_reg, col_reg}<16'b0000100011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000100011110000) && ({row_reg, col_reg}<16'b0000100011110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000100011110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100011110011) && ({row_reg, col_reg}<16'b0000100011110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100011110111) && ({row_reg, col_reg}<16'b0000100011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000100011111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100011111010) && ({row_reg, col_reg}<16'b0000100011111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000100011111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000100011111110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}==16'b0000100011111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100100000000) && ({row_reg, col_reg}<16'b0000100100000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100100000011) && ({row_reg, col_reg}<16'b0000100100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000100100001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100100001001) && ({row_reg, col_reg}<16'b0000100100001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100100001011) && ({row_reg, col_reg}<16'b0000100100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000100100001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100100001111) && ({row_reg, col_reg}<16'b0000100100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100100010010) && ({row_reg, col_reg}<16'b0000100100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000100100100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100100100110) && ({row_reg, col_reg}<16'b0000100100101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100100101010) && ({row_reg, col_reg}<16'b0000100100101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100100101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000100100101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100100101110) && ({row_reg, col_reg}<16'b0000100100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000100100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100100110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100100110010) && ({row_reg, col_reg}<16'b0000100100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100100110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000100100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100100110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000100100111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100100111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000100100111010) && ({row_reg, col_reg}<16'b0000100100111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100100111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000100100111101) && ({row_reg, col_reg}<16'b0000100100111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100100111111) && ({row_reg, col_reg}<16'b0000100101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100101000100) && ({row_reg, col_reg}<16'b0000100101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100101000111) && ({row_reg, col_reg}<16'b0000100101001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000100101001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000100101001010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000100101001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100101001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000100101001101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0000100101001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100101001111) && ({row_reg, col_reg}<16'b0000100101010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000100101010111) && ({row_reg, col_reg}<16'b0000100101011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100101011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000100101011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100101011011) && ({row_reg, col_reg}<16'b0000100101011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100101011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000100101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100101011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000100101100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100101100001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000100101100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000100101100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000100101100100) && ({row_reg, col_reg}<16'b0000100101101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100101101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000100101101001) && ({row_reg, col_reg}<16'b0000100101101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100101101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000100101101100) && ({row_reg, col_reg}<16'b0000100101110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000100101110001) && ({row_reg, col_reg}<16'b0000100101111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000100101111011) && ({row_reg, col_reg}<16'b0000100101111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100101111101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0000100101111110) && ({row_reg, col_reg}<16'b0000100110000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100110000000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000100110000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100110000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100110000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100110000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100110000101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000100110000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100110000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000100110001000) && ({row_reg, col_reg}<16'b0000100110001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100110001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000100110001101) && ({row_reg, col_reg}<16'b0000100110001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100110001111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000100110010000) && ({row_reg, col_reg}<16'b0000100110010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000100110010010) && ({row_reg, col_reg}<16'b0000100110010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000100110010101) && ({row_reg, col_reg}<16'b0000100110010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000100110010111) && ({row_reg, col_reg}<16'b0000100110011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100110011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000100110011101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000100110011110) && ({row_reg, col_reg}<16'b0000100110100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000100110100011) && ({row_reg, col_reg}<16'b0000100110100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000100110100111) && ({row_reg, col_reg}<16'b0000100110101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000100110101100) && ({row_reg, col_reg}<16'b0000100110110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000100110110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000100110110001) && ({row_reg, col_reg}<16'b0000100110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100110110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000100110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000100110110110) && ({row_reg, col_reg}<16'b0000100110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000100110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100110111001) && ({row_reg, col_reg}<16'b0000100110111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000100110111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000100110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100110111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000100110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000100111000000) && ({row_reg, col_reg}<16'b0000100111000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100111000010) && ({row_reg, col_reg}<16'b0000100111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000100111000100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000100111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100111000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000100111000111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000100111001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000100111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100111001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000100111001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000100111001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000100111001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000100111001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100111001111) && ({row_reg, col_reg}<16'b0000100111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100111010001) && ({row_reg, col_reg}<16'b0000100111110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000100111110000) && ({row_reg, col_reg}<16'b0000100111110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100111110011) && ({row_reg, col_reg}<16'b0000100111110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100111110111) && ({row_reg, col_reg}<16'b0000100111111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100111111001) && ({row_reg, col_reg}<16'b0000100111111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0000100111111011) && ({row_reg, col_reg}<16'b0000101000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101000000000) && ({row_reg, col_reg}<16'b0000101000000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000101000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101000000110) && ({row_reg, col_reg}<16'b0000101000001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000101000001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101000001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101000001011) && ({row_reg, col_reg}<16'b0000101000001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000101000001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101000001111) && ({row_reg, col_reg}<16'b0000101000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101000010010) && ({row_reg, col_reg}<16'b0000101000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000101000100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101000100110) && ({row_reg, col_reg}<16'b0000101000101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101000101110) && ({row_reg, col_reg}<16'b0000101000110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000101000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101000110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101000110010) && ({row_reg, col_reg}<16'b0000101000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101000110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000101000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101000110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000101000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101000111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000101000111010) && ({row_reg, col_reg}<16'b0000101000111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101000111100) && ({row_reg, col_reg}<16'b0000101001000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000101001000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000101001000100) && ({row_reg, col_reg}<16'b0000101001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101001000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000101001000111) && ({row_reg, col_reg}<16'b0000101001001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000101001001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101001001010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101001001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101001001100) && ({row_reg, col_reg}<16'b0000101001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000101001001111) && ({row_reg, col_reg}<16'b0000101001010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101001010111) && ({row_reg, col_reg}<16'b0000101001011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000101001011010) && ({row_reg, col_reg}<16'b0000101001011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101001011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000101001011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101001011111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000101001100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101001100001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000101001100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000101001100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000101001100100) && ({row_reg, col_reg}<16'b0000101001101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101001101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000101001101001) && ({row_reg, col_reg}<16'b0000101001101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101001101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101001101100) && ({row_reg, col_reg}<16'b0000101001101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101001101111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000101001110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000101001110001) && ({row_reg, col_reg}<16'b0000101001111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101001111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000101001111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000101001111101) && ({row_reg, col_reg}<16'b0000101010000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101010000000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000101010000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101010000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101010000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000101010000100) && ({row_reg, col_reg}<16'b0000101010000110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000101010000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101010000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000101010001000) && ({row_reg, col_reg}<16'b0000101010001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101010001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101010001110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000101010001111) && ({row_reg, col_reg}<16'b0000101010010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101010010010) && ({row_reg, col_reg}<16'b0000101010010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101010010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000101010010111) && ({row_reg, col_reg}<16'b0000101010011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101010011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101010011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000101010011101) && ({row_reg, col_reg}<16'b0000101010100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101010100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000101010100001) && ({row_reg, col_reg}<16'b0000101010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101010100011) && ({row_reg, col_reg}<16'b0000101010100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000101010100111) && ({row_reg, col_reg}<16'b0000101010101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101010101100) && ({row_reg, col_reg}<16'b0000101010110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000101010110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101010110001) && ({row_reg, col_reg}<16'b0000101010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101010110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000101010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000101010110110) && ({row_reg, col_reg}<16'b0000101010111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000101010111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000101010111101) && ({row_reg, col_reg}<16'b0000101011000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000101011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101011000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101011000010) && ({row_reg, col_reg}<16'b0000101011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000101011000100) && ({row_reg, col_reg}<16'b0000101011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000101011000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101011000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000101011001000) && ({row_reg, col_reg}<16'b0000101011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101011001010) && ({row_reg, col_reg}<16'b0000101011001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101011001111) && ({row_reg, col_reg}<16'b0000101011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101011010001) && ({row_reg, col_reg}<16'b0000101011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000101011110000) && ({row_reg, col_reg}<16'b0000101011110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000101011110011) && ({row_reg, col_reg}<16'b0000101011110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101011110111) && ({row_reg, col_reg}<16'b0000101011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000101011111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101011111010) && ({row_reg, col_reg}<16'b0000101011111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101011111110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}==16'b0000101011111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101100000000) && ({row_reg, col_reg}<16'b0000101100000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000101100000100) && ({row_reg, col_reg}<16'b0000101100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101100000110) && ({row_reg, col_reg}<16'b0000101100001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000101100001001) && ({row_reg, col_reg}<16'b0000101100001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101100001011) && ({row_reg, col_reg}<16'b0000101100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000101100001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101100001111) && ({row_reg, col_reg}<16'b0000101100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101100010010) && ({row_reg, col_reg}<16'b0000101100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000101100100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101100100110) && ({row_reg, col_reg}<16'b0000101100101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101100101110) && ({row_reg, col_reg}<16'b0000101100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000101100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101100110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101100110010) && ({row_reg, col_reg}<16'b0000101100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101100110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000101100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101100110111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000101100111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101100111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000101100111010) && ({row_reg, col_reg}<16'b0000101100111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101100111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000101100111101) && ({row_reg, col_reg}<16'b0000101100111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101100111111) && ({row_reg, col_reg}<16'b0000101101000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000101101000010) && ({row_reg, col_reg}<16'b0000101101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000101101000100) && ({row_reg, col_reg}<16'b0000101101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101101000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000101101000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101101001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000101101001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101101001010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000101101001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101101001100) && ({row_reg, col_reg}<16'b0000101101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000101101001111) && ({row_reg, col_reg}<16'b0000101101010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101101010101) && ({row_reg, col_reg}<16'b0000101101011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000101101011000) && ({row_reg, col_reg}<16'b0000101101011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101101011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101101011111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000101101100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101101100001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000101101100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000101101100011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0000101101100100) && ({row_reg, col_reg}<16'b0000101101101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101101101000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000101101101001) && ({row_reg, col_reg}<16'b0000101101101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101101101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101101101100) && ({row_reg, col_reg}<16'b0000101101110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000101101110001) && ({row_reg, col_reg}<16'b0000101101110100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101101110100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000101101110101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000101101110110)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0000101101110111) && ({row_reg, col_reg}<16'b0000101101111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101101111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000101101111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101101111101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000101101111110) && ({row_reg, col_reg}<16'b0000101110000000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000101110000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101110000001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000101110000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101110000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000101110000100) && ({row_reg, col_reg}<16'b0000101110000110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000101110000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101110000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101110001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101110001001) && ({row_reg, col_reg}<16'b0000101110001011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000101110001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101110001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101110001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101110001110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000101110001111) && ({row_reg, col_reg}<16'b0000101110010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101110010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000101110010010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000101110010011) && ({row_reg, col_reg}<16'b0000101110010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000101110010101) && ({row_reg, col_reg}<16'b0000101110010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000101110010111) && ({row_reg, col_reg}<16'b0000101110011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101110011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101110011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000101110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000101110011101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000101110011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101110011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101110100000) && ({row_reg, col_reg}<16'b0000101110100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000101110100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101110100011) && ({row_reg, col_reg}<16'b0000101110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000101110100110) && ({row_reg, col_reg}<16'b0000101110101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000101110101001) && ({row_reg, col_reg}<16'b0000101110101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101110101011) && ({row_reg, col_reg}<16'b0000101110110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000101110110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101110110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101110110010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000101110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101110110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000101110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000101110110110) && ({row_reg, col_reg}<16'b0000101110111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000101110111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101110111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000101110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000101110111111) && ({row_reg, col_reg}<16'b0000101111000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000101111000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101111000010) && ({row_reg, col_reg}<16'b0000101111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000101111000100) && ({row_reg, col_reg}<16'b0000101111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101111000110) && ({row_reg, col_reg}<16'b0000101111001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101111001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101111001011) && ({row_reg, col_reg}<16'b0000101111001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101111001101) && ({row_reg, col_reg}<16'b0000101111001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101111001111) && ({row_reg, col_reg}<16'b0000101111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101111010001) && ({row_reg, col_reg}<16'b0000101111101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000101111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101111110000) && ({row_reg, col_reg}<16'b0000101111110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000101111110011) && ({row_reg, col_reg}<16'b0000101111110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101111110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101111110110) && ({row_reg, col_reg}<16'b0000101111111010)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0000101111111010) && ({row_reg, col_reg}<16'b0000110000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110000000000) && ({row_reg, col_reg}<16'b0000110000000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000110000000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110000001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000110000001001) && ({row_reg, col_reg}<16'b0000110000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000110000001100) && ({row_reg, col_reg}<16'b0000110000001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000110000001110) && ({row_reg, col_reg}<16'b0000110000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110000010010) && ({row_reg, col_reg}<16'b0000110000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000110000100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110000100110) && ({row_reg, col_reg}<16'b0000110000101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110000101110) && ({row_reg, col_reg}<16'b0000110000110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000110000110000) && ({row_reg, col_reg}<16'b0000110000110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110000110010) && ({row_reg, col_reg}<16'b0000110000110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000110000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110000110111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000110000111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000110000111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000110000111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000110000111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110000111100) && ({row_reg, col_reg}<16'b0000110000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000110000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110000111111) && ({row_reg, col_reg}<16'b0000110001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000110001000001) && ({row_reg, col_reg}<16'b0000110001000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000110001000011) && ({row_reg, col_reg}<16'b0000110001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110001000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000110001000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110001001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000110001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110001001010) && ({row_reg, col_reg}<16'b0000110001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000110001001100) && ({row_reg, col_reg}<16'b0000110001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110001001111) && ({row_reg, col_reg}<16'b0000110001010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000110001010101) && ({row_reg, col_reg}<16'b0000110001011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110001011000) && ({row_reg, col_reg}<16'b0000110001011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110001011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110001011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110001011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000110001100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110001100001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000110001100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000110001100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110001100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000110001100101) && ({row_reg, col_reg}<16'b0000110001100111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000110001100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110001101000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0000110001101001) && ({row_reg, col_reg}<16'b0000110001101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110001101011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000110001101100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000110001101101) && ({row_reg, col_reg}<16'b0000110001110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110001110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000110001110001) && ({row_reg, col_reg}<16'b0000110001110100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110001110100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000110001110101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000110001110110)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000110001110111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110001111000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0000110001111001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0000110001111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110001111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000110001111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110001111101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000110001111110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000110001111111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000110010000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110010000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110010000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110010000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110010000100)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0000110010000101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000110010000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110010000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110010001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110010001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110010001010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000110010001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110010001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110010001110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000110010001111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000110010010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000110010010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000110010010010) && ({row_reg, col_reg}<16'b0000110010010100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000110010010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110010010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000110010010110) && ({row_reg, col_reg}<16'b0000110010011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110010011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000110010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000110010011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000110010011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000110010011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000110010100000) && ({row_reg, col_reg}<16'b0000110010100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000110010100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000110010100011) && ({row_reg, col_reg}<16'b0000110010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000110010100110) && ({row_reg, col_reg}<16'b0000110010101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110010101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000110010101010) && ({row_reg, col_reg}<16'b0000110010110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000110010110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110010110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110010110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000110010110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0000110010110100) && ({row_reg, col_reg}<16'b0000110010110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000110010110110) && ({row_reg, col_reg}<16'b0000110010111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000110010111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110010111010) && ({row_reg, col_reg}<16'b0000110010111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0000110010111100) && ({row_reg, col_reg}<16'b0000110010111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000110010111110) && ({row_reg, col_reg}<16'b0000110011000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110011000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000110011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110011000010) && ({row_reg, col_reg}<16'b0000110011000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110011000101) && ({row_reg, col_reg}<16'b0000110011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110011001111) && ({row_reg, col_reg}<16'b0000110011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110011010001) && ({row_reg, col_reg}<16'b0000110011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000110011101111) && ({row_reg, col_reg}<16'b0000110011110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000110011110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110011110100) && ({row_reg, col_reg}<16'b0000110011110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110011110110) && ({row_reg, col_reg}<16'b0000110011111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000110011111010) && ({row_reg, col_reg}<16'b0000110011111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110011111100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0000110011111101) && ({row_reg, col_reg}<16'b0000110100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110100000000) && ({row_reg, col_reg}<16'b0000110100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000110100001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110100001001) && ({row_reg, col_reg}<16'b0000110100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000110100001101) && ({row_reg, col_reg}<16'b0000110100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000110100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110100010010) && ({row_reg, col_reg}<16'b0000110100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000110100100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110100100110) && ({row_reg, col_reg}<16'b0000110100101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000110100101001) && ({row_reg, col_reg}<16'b0000110100101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110100101110) && ({row_reg, col_reg}<16'b0000110100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000110100110000) && ({row_reg, col_reg}<16'b0000110100110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110100110010) && ({row_reg, col_reg}<16'b0000110100110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000110100110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000110100110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000110100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110100110111) && ({row_reg, col_reg}<16'b0000110100111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000110100111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000110100111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000110100111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110100111100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0000110100111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000110100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110100111111) && ({row_reg, col_reg}<16'b0000110101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000110101000001) && ({row_reg, col_reg}<16'b0000110101000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000110101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110101000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000110101000111) && ({row_reg, col_reg}<16'b0000110101001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000110101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110101001010) && ({row_reg, col_reg}<16'b0000110101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000110101001100) && ({row_reg, col_reg}<16'b0000110101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110101001111) && ({row_reg, col_reg}<16'b0000110101010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000110101010101) && ({row_reg, col_reg}<16'b0000110101011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110101011000) && ({row_reg, col_reg}<16'b0000110101011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110101011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000110101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110101011111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000110101100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110101100001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000110101100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000110101100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000110101100100) && ({row_reg, col_reg}<16'b0000110101101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110101101000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0000110101101001) && ({row_reg, col_reg}<16'b0000110101101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110101101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000110101101100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000110101101101) && ({row_reg, col_reg}<16'b0000110101110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000110101110001) && ({row_reg, col_reg}<16'b0000110101110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000110101110101) && ({row_reg, col_reg}<16'b0000110101110111)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000110101110111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110101111000)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0000110101111001)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}>=16'b0000110101111010) && ({row_reg, col_reg}<16'b0000110101111100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0000110101111100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000110101111101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110101111110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000110101111111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000110110000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110110000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110110000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110110000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110110000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110110000101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000110110000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110110000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110110001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110110001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110110001010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000110110001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110110001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110110001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110110001110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000110110001111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000110110010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000110110010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000110110010010) && ({row_reg, col_reg}<16'b0000110110010100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000110110010100) && ({row_reg, col_reg}<16'b0000110110010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110110010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000110110010111) && ({row_reg, col_reg}<16'b0000110110011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110110011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110110011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110110011100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000110110011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000110110011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000110110011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000110110100000) && ({row_reg, col_reg}<16'b0000110110100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000110110100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000110110100011) && ({row_reg, col_reg}<16'b0000110110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000110110100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0000110110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110110101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110110101010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000110110101011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000110110101100) && ({row_reg, col_reg}<16'b0000110110101110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000110110101110) && ({row_reg, col_reg}<16'b0000110110110000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000110110110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110110110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110110110010)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0000110110110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0000110110110100) && ({row_reg, col_reg}<16'b0000110110110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000110110110110) && ({row_reg, col_reg}<16'b0000110110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0000110110111000) && ({row_reg, col_reg}<16'b0000110110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110110111010) && ({row_reg, col_reg}<16'b0000110110111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0000110110111100) && ({row_reg, col_reg}<16'b0000110111000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000110111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110111000010) && ({row_reg, col_reg}<16'b0000110111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110111000110) && ({row_reg, col_reg}<16'b0000110111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110111001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000110111001111) && ({row_reg, col_reg}<16'b0000110111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110111010001) && ({row_reg, col_reg}<16'b0000110111101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000110111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110111110000) && ({row_reg, col_reg}<16'b0000110111110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000110111110010) && ({row_reg, col_reg}<16'b0000110111110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110111110111) && ({row_reg, col_reg}<16'b0000110111111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000110111111010) && ({row_reg, col_reg}<16'b0000110111111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110111111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000110111111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110111111110)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}==16'b0000110111111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111000000000) && ({row_reg, col_reg}<16'b0000111000001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000111000001001) && ({row_reg, col_reg}<16'b0000111000001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000111000001111) && ({row_reg, col_reg}<16'b0000111000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000111000100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000111000100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111000100111) && ({row_reg, col_reg}<16'b0000111000101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000111000101001) && ({row_reg, col_reg}<16'b0000111000101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111000101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000111000101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111000101110) && ({row_reg, col_reg}<16'b0000111000110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000111000110000) && ({row_reg, col_reg}<16'b0000111000110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111000110010) && ({row_reg, col_reg}<16'b0000111000110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111000110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111000110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000111000111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111000111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000111000111010) && ({row_reg, col_reg}<16'b0000111000111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111000111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111000111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000111000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111000111111) && ({row_reg, col_reg}<16'b0000111001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000111001000001) && ({row_reg, col_reg}<16'b0000111001000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111001000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000111001000100) && ({row_reg, col_reg}<16'b0000111001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111001000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000111001000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111001001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000111001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000111001001010) && ({row_reg, col_reg}<16'b0000111001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000111001001100) && ({row_reg, col_reg}<16'b0000111001001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000111001001111) && ({row_reg, col_reg}<16'b0000111001010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000111001010110) && ({row_reg, col_reg}<16'b0000111001011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111001011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000111001011001) && ({row_reg, col_reg}<16'b0000111001011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000111001011011) && ({row_reg, col_reg}<16'b0000111001011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111001011101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000111001011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111001011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000111001100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111001100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111001100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000111001100011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0000111001100100) && ({row_reg, col_reg}<16'b0000111001100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111001100111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000111001101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000111001101001) && ({row_reg, col_reg}<16'b0000111001101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111001101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000111001101100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000111001101101) && ({row_reg, col_reg}<16'b0000111001110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111001110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000111001110001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000111001110010) && ({row_reg, col_reg}<16'b0000111001110100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111001110100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000111001110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000111001110110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000111001110111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000111001111000) && ({row_reg, col_reg}<16'b0000111001111011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0000111001111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111001111100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000111001111101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111001111110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000111001111111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000111010000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111010000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111010000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000111010000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111010000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111010000101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000111010000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111010000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111010001000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000111010001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111010001010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000111010001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111010001101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000111010001110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111010001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111010010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000111010010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111010010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111010010011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000111010010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111010010101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0000111010010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000111010010111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000111010011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111010011001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000111010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000111010011011) && ({row_reg, col_reg}<16'b0000111010011101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111010011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111010011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111010011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000111010100000) && ({row_reg, col_reg}<16'b0000111010100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000111010100010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0000111010100011) && ({row_reg, col_reg}<16'b0000111010100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000111010100101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0000111010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000111010100111) && ({row_reg, col_reg}<16'b0000111010110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111010110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000111010110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111010110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0000111010111000) && ({row_reg, col_reg}<16'b0000111010111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111010111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000111010111101) && ({row_reg, col_reg}<16'b0000111010111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000111010111111) && ({row_reg, col_reg}<16'b0000111011000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000111011000001) && ({row_reg, col_reg}<16'b0000111011000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111011000011) && ({row_reg, col_reg}<16'b0000111011000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111011000101) && ({row_reg, col_reg}<16'b0000111011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111011010001) && ({row_reg, col_reg}<16'b0000111011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000111011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000111011110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111011110100) && ({row_reg, col_reg}<16'b0000111011111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111011111000) && ({row_reg, col_reg}<16'b0000111011111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000111011111010) && ({row_reg, col_reg}<16'b0000111011111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111011111110)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}==16'b0000111011111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111100000000) && ({row_reg, col_reg}<16'b0000111100001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000111100001010) && ({row_reg, col_reg}<16'b0000111100001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111100001100) && ({row_reg, col_reg}<16'b0000111100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111100010001) && ({row_reg, col_reg}<16'b0000111100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000111100100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111100100110) && ({row_reg, col_reg}<16'b0000111100101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000111100101001) && ({row_reg, col_reg}<16'b0000111100101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111100101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000111100101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111100101110) && ({row_reg, col_reg}<16'b0000111100110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000111100110000) && ({row_reg, col_reg}<16'b0000111100110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111100110010) && ({row_reg, col_reg}<16'b0000111100110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111100110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111100110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111100111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111100111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111100111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111100111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111100111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000111100111110) && ({row_reg, col_reg}<16'b0000111101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111101000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000111101000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111101000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000111101000100) && ({row_reg, col_reg}<16'b0000111101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111101000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111101001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111101001011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0000111101001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111101001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111101001110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000111101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000111101010000) && ({row_reg, col_reg}<16'b0000111101011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000111101011000) && ({row_reg, col_reg}<16'b0000111101011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000111101011100) && ({row_reg, col_reg}<16'b0000111101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111101011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000111101011111) && ({row_reg, col_reg}<16'b0000111101100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111101100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111101100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000111101100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000111101100100) && ({row_reg, col_reg}<16'b0000111101100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111101100111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000111101101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000111101101001) && ({row_reg, col_reg}<16'b0000111101101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111101101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111101101101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000111101101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000111101101111) && ({row_reg, col_reg}<16'b0000111101110001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000111101110001) && ({row_reg, col_reg}<16'b0000111101111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000111101111001) && ({row_reg, col_reg}<16'b0000111101111100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111101111100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000111101111101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111101111110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000111101111111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000111110000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111110000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111110000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000111110000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111110000100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000111110000101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000111110000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000111110000111) && ({row_reg, col_reg}<16'b0000111110001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111110001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111110001100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000111110001101) && ({row_reg, col_reg}<16'b0000111110001111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000111110001111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000111110010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000111110010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111110010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111110010011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000111110010100) && ({row_reg, col_reg}<16'b0000111110010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000111110010110) && ({row_reg, col_reg}<16'b0000111110011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000111110011000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0000111110011001) && ({row_reg, col_reg}<16'b0000111110011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111110011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000111110011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111110011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000111110011110) && ({row_reg, col_reg}<16'b0000111110100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000111110100000) && ({row_reg, col_reg}<16'b0000111110100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000111110100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000111110100011) && ({row_reg, col_reg}<16'b0000111110100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000111110100111) && ({row_reg, col_reg}<16'b0000111110110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111110110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000111110110110) && ({row_reg, col_reg}<16'b0000111110111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111110111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000111110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000111110111011) && ({row_reg, col_reg}<16'b0000111110111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000111110111101) && ({row_reg, col_reg}<16'b0000111111000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111111000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000111111000001) && ({row_reg, col_reg}<16'b0000111111000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111111000110) && ({row_reg, col_reg}<16'b0000111111001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000111111001000) && ({row_reg, col_reg}<16'b0000111111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111111010001) && ({row_reg, col_reg}<16'b0000111111101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000111111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111111110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111111110010) && ({row_reg, col_reg}<16'b0000111111110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000111111110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111111110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111111110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000111111110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111111111000) && ({row_reg, col_reg}<16'b0000111111111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000111111111010) && ({row_reg, col_reg}<16'b0000111111111101)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0000111111111101) && ({row_reg, col_reg}<16'b0001000000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000000000000) && ({row_reg, col_reg}<16'b0001000000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000000000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001000000000111) && ({row_reg, col_reg}<16'b0001000000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000000001101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001000000001110) && ({row_reg, col_reg}<16'b0001000000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000000010010) && ({row_reg, col_reg}<16'b0001000000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001000000100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000000100110) && ({row_reg, col_reg}<16'b0001000000101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000000101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000000101001) && ({row_reg, col_reg}<16'b0001000000101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000000101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000000101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001000000110000) && ({row_reg, col_reg}<16'b0001000000110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000000110010) && ({row_reg, col_reg}<16'b0001000000110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000000110100) && ({row_reg, col_reg}<16'b0001000000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001000000110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000000110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000000111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000000111001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0001000000111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000000111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000000111100)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b0001000000111101) && ({row_reg, col_reg}<16'b0001000001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000001000001) && ({row_reg, col_reg}<16'b0001000001000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001000001000100) && ({row_reg, col_reg}<16'b0001000001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000001000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000001000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000001001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001000001001001) && ({row_reg, col_reg}<16'b0001000001001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000001001100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001000001001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000001001110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001000001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001000001010000) && ({row_reg, col_reg}<16'b0001000001010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001000001010111) && ({row_reg, col_reg}<16'b0001000001011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000001011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000001011101)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0001000001011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001000001011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000001100000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001000001100001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001000001100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001000001100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001000001100100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001000001100101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001000001100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000001100111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001000001101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001000001101001) && ({row_reg, col_reg}<16'b0001000001101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000001101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000001101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000001101110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001000001101111) && ({row_reg, col_reg}<16'b0001000001110001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001000001110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000001110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001000001110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001000001110100) && ({row_reg, col_reg}<16'b0001000001110110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001000001110110) && ({row_reg, col_reg}<16'b0001000001111000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000001111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001000001111001) && ({row_reg, col_reg}<16'b0001000001111011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001000001111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001000001111100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001000001111101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001000001111110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001000001111111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001000010000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001000010000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000010000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001000010000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000010000100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001000010000101)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0001000010000110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001000010000111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001000010001000) && ({row_reg, col_reg}<16'b0001000010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000010001100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001000010001101) && ({row_reg, col_reg}<16'b0001000010001111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001000010001111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001000010010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001000010010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000010010010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001000010010011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001000010010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001000010010101) && ({row_reg, col_reg}<16'b0001000010011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001000010011000) && ({row_reg, col_reg}<16'b0001000010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000010011010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001000010011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001000010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001000010011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000010011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000010011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001000010100000) && ({row_reg, col_reg}<16'b0001000010100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001000010100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001000010100011) && ({row_reg, col_reg}<16'b0001000010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001000010100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0001000010100111) && ({row_reg, col_reg}<16'b0001000010101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001000010101100) && ({row_reg, col_reg}<16'b0001000010110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001000010110010) && ({row_reg, col_reg}<16'b0001000010110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000010110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001000010110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000010110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001000010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000010111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001000010111010) && ({row_reg, col_reg}<16'b0001000010111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001000010111100) && ({row_reg, col_reg}<16'b0001000010111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001000010111110) && ({row_reg, col_reg}<16'b0001000011000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001000011000000) && ({row_reg, col_reg}<16'b0001000011000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000011000010) && ({row_reg, col_reg}<16'b0001000011000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000011000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000011000111) && ({row_reg, col_reg}<16'b0001000011001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001000011001001) && ({row_reg, col_reg}<16'b0001000011001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000011001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000011001100) && ({row_reg, col_reg}<16'b0001000011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000011010001) && ({row_reg, col_reg}<16'b0001000011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001000011101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001000011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001000011110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000011110100) && ({row_reg, col_reg}<16'b0001000011111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000011111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000011111001) && ({row_reg, col_reg}<16'b0001000011111100)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0001000011111100) && ({row_reg, col_reg}<16'b0001000100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000100000000) && ({row_reg, col_reg}<16'b0001000100000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000100000010) && ({row_reg, col_reg}<16'b0001000100000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000100000100) && ({row_reg, col_reg}<16'b0001000100001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000100001110) && ({row_reg, col_reg}<16'b0001000100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000100010011) && ({row_reg, col_reg}<16'b0001000100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001000100100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000100100110) && ({row_reg, col_reg}<16'b0001000100101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000100101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000100101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001000100101011) && ({row_reg, col_reg}<16'b0001000100101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000100101110) && ({row_reg, col_reg}<16'b0001000100110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000100110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000100110010) && ({row_reg, col_reg}<16'b0001000100110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000100110100) && ({row_reg, col_reg}<16'b0001000100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001000100110110) && ({row_reg, col_reg}<16'b0001000100111000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001000100111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000100111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000100111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000100111011) && ({row_reg, col_reg}<16'b0001000101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000101000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001000101000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000101000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001000101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000101000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000101001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001000101001001) && ({row_reg, col_reg}<16'b0001000101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000101001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001000101001100)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==16'b0001000101001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000101001110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001000101001111) && ({row_reg, col_reg}<16'b0001000101010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000101010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001000101010110) && ({row_reg, col_reg}<16'b0001000101011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001000101011000) && ({row_reg, col_reg}<16'b0001000101011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000101011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001000101011101) && ({row_reg, col_reg}<16'b0001000101011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001000101011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000101100000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001000101100001) && ({row_reg, col_reg}<16'b0001000101100011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001000101100011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001000101100100) && ({row_reg, col_reg}<16'b0001000101100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001000101100110) && ({row_reg, col_reg}<16'b0001000101101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000101101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001000101101001) && ({row_reg, col_reg}<16'b0001000101101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000101101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000101101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001000101101101) && ({row_reg, col_reg}<16'b0001000101101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001000101101111) && ({row_reg, col_reg}<16'b0001000101110001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001000101110001)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0001000101110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001000101110011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001000101110100) && ({row_reg, col_reg}<16'b0001000101110110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001000101110110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001000101110111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001000101111000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001000101111001)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0001000101111010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001000101111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001000101111100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001000101111101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001000101111110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001000101111111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001000110000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001000110000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000110000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001000110000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000110000100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001000110000101)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0001000110000110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001000110000111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001000110001000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001000110001001) && ({row_reg, col_reg}<16'b0001000110001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000110001011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001000110001100) && ({row_reg, col_reg}<16'b0001000110001111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001000110001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001000110010000) && ({row_reg, col_reg}<16'b0001000110010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001000110010010) && ({row_reg, col_reg}<16'b0001000110010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001000110010101) && ({row_reg, col_reg}<16'b0001000110011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001000110011000) && ({row_reg, col_reg}<16'b0001000110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001000110011010) && ({row_reg, col_reg}<16'b0001000110011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001000110011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000110011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000110011110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001000110011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000110100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001000110100001) && ({row_reg, col_reg}<16'b0001000110100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000110100011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0001000110100100) && ({row_reg, col_reg}<16'b0001000110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001000110100110) && ({row_reg, col_reg}<16'b0001000110101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001000110101100) && ({row_reg, col_reg}<16'b0001000110101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000110101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001000110101111) && ({row_reg, col_reg}<16'b0001000110110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000110110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001000110110011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0001000110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001000110110110) && ({row_reg, col_reg}<16'b0001000110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001000110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000110111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001000110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001000110111011) && ({row_reg, col_reg}<16'b0001000110111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001000110111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000110111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001000111000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001000111000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000111000010) && ({row_reg, col_reg}<16'b0001000111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000111000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000111000110) && ({row_reg, col_reg}<16'b0001000111001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001000111001000) && ({row_reg, col_reg}<16'b0001000111001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000111001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000111001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000111001100) && ({row_reg, col_reg}<16'b0001000111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000111001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000111001111) && ({row_reg, col_reg}<16'b0001000111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000111010001) && ({row_reg, col_reg}<16'b0001000111101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001000111101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001000111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000111110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000111110010) && ({row_reg, col_reg}<16'b0001000111110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000111110100) && ({row_reg, col_reg}<16'b0001000111110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000111110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000111111000) && ({row_reg, col_reg}<16'b0001000111111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000111111101)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0001000111111110) && ({row_reg, col_reg}<16'b0001001000000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001000000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001001000000011) && ({row_reg, col_reg}<16'b0001001000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001000000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001000000110) && ({row_reg, col_reg}<16'b0001001000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001000001111) && ({row_reg, col_reg}<16'b0001001000010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001000010011) && ({row_reg, col_reg}<16'b0001001000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001001000100101) && ({row_reg, col_reg}<16'b0001001000100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001000100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001000101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001000101001) && ({row_reg, col_reg}<16'b0001001000101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001000101011) && ({row_reg, col_reg}<16'b0001001000101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001000101110) && ({row_reg, col_reg}<16'b0001001000110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001000110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001000110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001000110100) && ({row_reg, col_reg}<16'b0001001000111000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001001000111000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0001001000111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001000111010) && ({row_reg, col_reg}<16'b0001001000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001000111110) && ({row_reg, col_reg}<16'b0001001001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001001000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001001001000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001001000011) && ({row_reg, col_reg}<16'b0001001001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001001000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001001000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001001001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001001001100) && ({row_reg, col_reg}<16'b0001001001001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001001001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001001010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001001001010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001001010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001001001010011) && ({row_reg, col_reg}<16'b0001001001010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001001010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001001010110) && ({row_reg, col_reg}<16'b0001001001011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001001001011101) && ({row_reg, col_reg}<16'b0001001001011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001001001011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001001001100000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001001001100001) && ({row_reg, col_reg}<16'b0001001001100011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001001001100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001001001100100) && ({row_reg, col_reg}<16'b0001001001100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001001100110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001001001100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001001001101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001001001101001) && ({row_reg, col_reg}<16'b0001001001101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001001101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001001001101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001001001101101) && ({row_reg, col_reg}<16'b0001001001101111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001001001101111) && ({row_reg, col_reg}<16'b0001001001110001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001001001110001)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0001001001110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001001001110011) && ({row_reg, col_reg}<16'b0001001001111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001001001111000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001001001111001)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0001001001111010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001001001111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001001001111100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001001001111101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001001001111110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001001001111111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001001010000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001001010000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001001010000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001001010000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001001010000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001001010000101) && ({row_reg, col_reg}<16'b0001001010000111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001001010000111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001001010001000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001001010001001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0001001010001010) && ({row_reg, col_reg}<16'b0001001010001100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001001010001100)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0001001010001101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0001001010001110)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0001001010001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001001010010000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0001001010010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001001010010010) && ({row_reg, col_reg}<16'b0001001010010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001001010010100) && ({row_reg, col_reg}<16'b0001001010011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001001010011000) && ({row_reg, col_reg}<16'b0001001010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001001010011010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001001010011011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001001010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001001010011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001010011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001010011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001010100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001001010100001) && ({row_reg, col_reg}<16'b0001001010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001010100011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0001001010100100) && ({row_reg, col_reg}<16'b0001001010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001001010100110) && ({row_reg, col_reg}<16'b0001001010110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001001010110000) && ({row_reg, col_reg}<16'b0001001010110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001010110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001001010110011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0001001010110100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0001001010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001001010110110) && ({row_reg, col_reg}<16'b0001001010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001001010111000) && ({row_reg, col_reg}<16'b0001001010111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001010111100) && ({row_reg, col_reg}<16'b0001001010111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001001010111110) && ({row_reg, col_reg}<16'b0001001011000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001011000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001001011000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001011000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001001011000100) && ({row_reg, col_reg}<16'b0001001011000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001011000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001001011000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001011001000) && ({row_reg, col_reg}<16'b0001001011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001001011001100) && ({row_reg, col_reg}<16'b0001001011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001001011001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001001011001111) && ({row_reg, col_reg}<16'b0001001011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001011010001) && ({row_reg, col_reg}<16'b0001001011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001001011101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001001011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001011110010) && ({row_reg, col_reg}<16'b0001001011110100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0001001011110100) && ({row_reg, col_reg}<16'b0001001100000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001001100000011) && ({row_reg, col_reg}<16'b0001001100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001100000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001100000111) && ({row_reg, col_reg}<16'b0001001100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001100010011) && ({row_reg, col_reg}<16'b0001001100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001001100100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001100100110) && ({row_reg, col_reg}<16'b0001001100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001001100101000) && ({row_reg, col_reg}<16'b0001001100101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001100101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001001100101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001100101110) && ({row_reg, col_reg}<16'b0001001100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001001100110000) && ({row_reg, col_reg}<16'b0001001100110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001100110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001100110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001100110100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001001100110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001001100110110) && ({row_reg, col_reg}<16'b0001001100111001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001001100111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001001100111010) && ({row_reg, col_reg}<16'b0001001100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001100111110) && ({row_reg, col_reg}<16'b0001001101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001101000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001001101000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001101000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001101000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001101000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001101000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001101001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001101001100) && ({row_reg, col_reg}<16'b0001001101001110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001001101001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001101001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001001101010000) && ({row_reg, col_reg}<16'b0001001101010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001001101010011) && ({row_reg, col_reg}<16'b0001001101011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001001101011101) && ({row_reg, col_reg}<16'b0001001101011111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001001101011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001001101100000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001001101100001) && ({row_reg, col_reg}<16'b0001001101100011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001001101100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001001101100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001001101100101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001001101100110) && ({row_reg, col_reg}<16'b0001001101101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001001101101000) && ({row_reg, col_reg}<16'b0001001101101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001101101010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0001001101101011) && ({row_reg, col_reg}<16'b0001001101101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001001101101101) && ({row_reg, col_reg}<16'b0001001101101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001001101101111) && ({row_reg, col_reg}<16'b0001001101110001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001001101110001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001001101110010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001001101110011) && ({row_reg, col_reg}<16'b0001001101111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001001101111000) && ({row_reg, col_reg}<16'b0001001101111011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001001101111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001001101111100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001001101111101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001001101111110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001001101111111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001001110000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001001110000001) && ({row_reg, col_reg}<16'b0001001110000011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001001110000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001001110000100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001001110000101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0001001110000110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0001001110000111) && ({row_reg, col_reg}<16'b0001001110001001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001001110001001)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0001001110001010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001001110001011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001001110001100)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0001001110001101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0001001110001110)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0001001110001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001001110010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001001110010001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001001110010010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001001110010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001001110010100) && ({row_reg, col_reg}<16'b0001001110011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001001110011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001001110011001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001001110011010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001001110011011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001001110011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001001110011101) && ({row_reg, col_reg}<16'b0001001110100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001110100000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001001110100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001001110100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001110100011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0001001110100100) && ({row_reg, col_reg}<16'b0001001110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001001110100110) && ({row_reg, col_reg}<16'b0001001110101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001001110101010) && ({row_reg, col_reg}<16'b0001001110101100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001001110101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001001110101101) && ({row_reg, col_reg}<16'b0001001110110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001001110110000) && ({row_reg, col_reg}<16'b0001001110110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001110110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001001110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001001110110110) && ({row_reg, col_reg}<16'b0001001110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001001110111000) && ({row_reg, col_reg}<16'b0001001110111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001110111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001001110111100) && ({row_reg, col_reg}<16'b0001001110111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001001110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001110111111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0001001111000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001111000001) && ({row_reg, col_reg}<16'b0001001111000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001111000011) && ({row_reg, col_reg}<16'b0001001111000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001001111000111) && ({row_reg, col_reg}<16'b0001001111001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001001111001001) && ({row_reg, col_reg}<16'b0001001111001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001111001011) && ({row_reg, col_reg}<16'b0001001111001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001111001111) && ({row_reg, col_reg}<16'b0001001111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001111010001) && ({row_reg, col_reg}<16'b0001001111101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001001111101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001001111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001111110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001111110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001111110011) && ({row_reg, col_reg}<16'b0001001111111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001111111100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0001001111111101) && ({row_reg, col_reg}<16'b0001010000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010000000110) && ({row_reg, col_reg}<16'b0001010000001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001010000001000) && ({row_reg, col_reg}<16'b0001010000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010000010011) && ({row_reg, col_reg}<16'b0001010000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001010000100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010000100110) && ({row_reg, col_reg}<16'b0001010000101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001010000101001) && ({row_reg, col_reg}<16'b0001010000101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010000101110) && ({row_reg, col_reg}<16'b0001010000110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001010000110000) && ({row_reg, col_reg}<16'b0001010000110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010000110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010000110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010000110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001010000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010000110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001010000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010000111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001010000111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010000111011) && ({row_reg, col_reg}<16'b0001010001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010001000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001010001000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001010001000011) && ({row_reg, col_reg}<16'b0001010001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010001000110) && ({row_reg, col_reg}<16'b0001010001001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001010001001001) && ({row_reg, col_reg}<16'b0001010001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001010001001100) && ({row_reg, col_reg}<16'b0001010001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010001001111) && ({row_reg, col_reg}<16'b0001010001010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001010001010001) && ({row_reg, col_reg}<16'b0001010001010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001010001010011) && ({row_reg, col_reg}<16'b0001010001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010001011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010001100000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001010001100001) && ({row_reg, col_reg}<16'b0001010001100011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001010001100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001010001100100) && ({row_reg, col_reg}<16'b0001010001100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010001100111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001010001101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001010001101001) && ({row_reg, col_reg}<16'b0001010001101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010001101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001010001101100) && ({row_reg, col_reg}<16'b0001010001101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001010001101111) && ({row_reg, col_reg}<16'b0001010001110011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001010001110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010001110100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001010001110101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0001010001110110) && ({row_reg, col_reg}<16'b0001010001111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001010001111000) && ({row_reg, col_reg}<16'b0001010001111011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001010001111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010001111100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001010001111101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010001111110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001010001111111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001010010000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001010010000001) && ({row_reg, col_reg}<16'b0001010010000011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001010010000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010010000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010010000101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0001010010000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010010000111)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0001010010001000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001010010001001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0001010010001010)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0001010010001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010010001100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001010010001101)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0001010010001110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001010010001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010010010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001010010010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010010010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010010010011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001010010010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001010010010101) && ({row_reg, col_reg}<16'b0001010010011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001010010011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010010011001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001010010011010) && ({row_reg, col_reg}<16'b0001010010011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001010010011101) && ({row_reg, col_reg}<16'b0001010010100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001010010100000) && ({row_reg, col_reg}<16'b0001010010100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001010010100010) && ({row_reg, col_reg}<16'b0001010010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001010010100110) && ({row_reg, col_reg}<16'b0001010010101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001010010101001) && ({row_reg, col_reg}<16'b0001010010101011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001010010101011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001010010101100) && ({row_reg, col_reg}<16'b0001010010110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010010110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001010010110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010010110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001010010110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001010010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001010010110110) && ({row_reg, col_reg}<16'b0001010010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001010010111000) && ({row_reg, col_reg}<16'b0001010010111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010010111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001010010111100) && ({row_reg, col_reg}<16'b0001010010111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001010010111110) && ({row_reg, col_reg}<16'b0001010011000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010011000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001010011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010011000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010011000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010011000100) && ({row_reg, col_reg}<16'b0001010011000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001010011000111) && ({row_reg, col_reg}<16'b0001010011001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001010011001001) && ({row_reg, col_reg}<16'b0001010011001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010011001101) && ({row_reg, col_reg}<16'b0001010011001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001010011001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010011010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010011010001) && ({row_reg, col_reg}<16'b0001010011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001010011101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001010011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001010011110001) && ({row_reg, col_reg}<16'b0001010011110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010011110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001010011111000) && ({row_reg, col_reg}<16'b0001010011111111)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}==16'b0001010011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001010100000000) && ({row_reg, col_reg}<16'b0001010100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010100000110) && ({row_reg, col_reg}<16'b0001010100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001010100001000) && ({row_reg, col_reg}<16'b0001010100001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010100001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001010100001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010100001100) && ({row_reg, col_reg}<16'b0001010100001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001010100001110) && ({row_reg, col_reg}<16'b0001010100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010100010011) && ({row_reg, col_reg}<16'b0001010100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001010100100101) && ({row_reg, col_reg}<16'b0001010100100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010100100111) && ({row_reg, col_reg}<16'b0001010100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001010100101001) && ({row_reg, col_reg}<16'b0001010100110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010100110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001010100110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010100110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001010100110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010100110111) && ({row_reg, col_reg}<16'b0001010100111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001010100111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001010100111010) && ({row_reg, col_reg}<16'b0001010101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001010101000001) && ({row_reg, col_reg}<16'b0001010101000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010101000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010101000100) && ({row_reg, col_reg}<16'b0001010101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010101000111) && ({row_reg, col_reg}<16'b0001010101001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001010101001001) && ({row_reg, col_reg}<16'b0001010101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010101001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010101001101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0001010101001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010101001111) && ({row_reg, col_reg}<16'b0001010101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010101011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001010101011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010101100000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001010101100001) && ({row_reg, col_reg}<16'b0001010101100011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001010101100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001010101100100) && ({row_reg, col_reg}<16'b0001010101100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010101100110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001010101100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010101101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001010101101001) && ({row_reg, col_reg}<16'b0001010101101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010101101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001010101101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010101101101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001010101101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010101101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001010101110000) && ({row_reg, col_reg}<16'b0001010101110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010101110011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0001010101110100) && ({row_reg, col_reg}<16'b0001010101110110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0001010101110110) && ({row_reg, col_reg}<16'b0001010101111000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0001010101111000) && ({row_reg, col_reg}<16'b0001010101111011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001010101111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010101111100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001010101111101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001010101111110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001010101111111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001010110000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001010110000001) && ({row_reg, col_reg}<16'b0001010110000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001010110000011) && ({row_reg, col_reg}<16'b0001010110000101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010110000101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0001010110000110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001010110000111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001010110001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001010110001001) && ({row_reg, col_reg}<16'b0001010110001011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001010110001011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001010110001100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010110001101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001010110001110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010110001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010110010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001010110010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001010110010010) && ({row_reg, col_reg}<16'b0001010110010100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010110010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001010110010101) && ({row_reg, col_reg}<16'b0001010110011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001010110011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010110011001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001010110011010) && ({row_reg, col_reg}<16'b0001010110011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001010110011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010110011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010110011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001010110100000) && ({row_reg, col_reg}<16'b0001010110100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001010110100011) && ({row_reg, col_reg}<16'b0001010110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001010110100110) && ({row_reg, col_reg}<16'b0001010110101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001010110101011) && ({row_reg, col_reg}<16'b0001010110110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010110110001)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0001010110110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001010110110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001010110110100) && ({row_reg, col_reg}<16'b0001010110110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010110110111) && ({row_reg, col_reg}<16'b0001010110111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001010110111100) && ({row_reg, col_reg}<16'b0001010111000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001010111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010111000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010111000011) && ({row_reg, col_reg}<16'b0001010111000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001010111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010111000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010111001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001010111001001) && ({row_reg, col_reg}<16'b0001010111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010111001110) && ({row_reg, col_reg}<16'b0001010111010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010111010001) && ({row_reg, col_reg}<16'b0001010111101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001010111101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001010111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010111110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001010111110001) && ({row_reg, col_reg}<16'b0001010111110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010111110111) && ({row_reg, col_reg}<16'b0001010111111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001010111111001) && ({row_reg, col_reg}<16'b0001010111111111)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}==16'b0001010111111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001011000000000) && ({row_reg, col_reg}<16'b0001011000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011000000101) && ({row_reg, col_reg}<16'b0001011000000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001011000000111) && ({row_reg, col_reg}<16'b0001011000001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011000001001) && ({row_reg, col_reg}<16'b0001011000001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011000001011) && ({row_reg, col_reg}<16'b0001011000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011000001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011000001110) && ({row_reg, col_reg}<16'b0001011000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011000010011) && ({row_reg, col_reg}<16'b0001011000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001011000100101) && ({row_reg, col_reg}<16'b0001011000101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011000101000) && ({row_reg, col_reg}<16'b0001011000101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011000101100) && ({row_reg, col_reg}<16'b0001011000110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011000110010) && ({row_reg, col_reg}<16'b0001011000110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001011000110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001011000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011000110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001011000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011000111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001011000111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011000111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001011000111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011000111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001011000111110) && ({row_reg, col_reg}<16'b0001011001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011001000001) && ({row_reg, col_reg}<16'b0001011001000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001011001000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011001000100) && ({row_reg, col_reg}<16'b0001011001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011001000111) && ({row_reg, col_reg}<16'b0001011001001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001011001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011001001010) && ({row_reg, col_reg}<16'b0001011001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011001001100) && ({row_reg, col_reg}<16'b0001011001010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011001010000) && ({row_reg, col_reg}<16'b0001011001011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011001011000) && ({row_reg, col_reg}<16'b0001011001011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011001011010) && ({row_reg, col_reg}<16'b0001011001011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011001011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001011001011111) && ({row_reg, col_reg}<16'b0001011001100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011001100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001011001100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001011001100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001011001100100) && ({row_reg, col_reg}<16'b0001011001100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011001100111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001011001101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001011001101001) && ({row_reg, col_reg}<16'b0001011001101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011001101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001011001101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011001101101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001011001101110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001011001101111) && ({row_reg, col_reg}<16'b0001011001110001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001011001110001) && ({row_reg, col_reg}<16'b0001011001111011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001011001111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001011001111100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001011001111101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001011001111110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001011001111111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001011010000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001011010000001) && ({row_reg, col_reg}<16'b0001011010000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011010000011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001011010000100) && ({row_reg, col_reg}<16'b0001011010000110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001011010000110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001011010000111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001011010001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011010001001) && ({row_reg, col_reg}<16'b0001011010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011010001100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001011010001101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001011010001110)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0001011010001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011010010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001011010010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001011010010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001011010010011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001011010010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001011010010101) && ({row_reg, col_reg}<16'b0001011010011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001011010011000) && ({row_reg, col_reg}<16'b0001011010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001011010011010) && ({row_reg, col_reg}<16'b0001011010011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001011010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001011010011101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001011010011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011010011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011010100000) && ({row_reg, col_reg}<16'b0001011010100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001011010100010) && ({row_reg, col_reg}<16'b0001011010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001011010100110) && ({row_reg, col_reg}<16'b0001011010101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011010101011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001011010101100) && ({row_reg, col_reg}<16'b0001011010110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001011010110001) && ({row_reg, col_reg}<16'b0001011010110011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001011010110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001011010110100) && ({row_reg, col_reg}<16'b0001011010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001011010111001) && ({row_reg, col_reg}<16'b0001011010111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011010111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001011010111100) && ({row_reg, col_reg}<16'b0001011011000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001011011000000) && ({row_reg, col_reg}<16'b0001011011000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011011000011) && ({row_reg, col_reg}<16'b0001011011000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001011011000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011011000110) && ({row_reg, col_reg}<16'b0001011011001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001011011001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001011011001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011011001010) && ({row_reg, col_reg}<16'b0001011011001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011011001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001011011001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011011001110) && ({row_reg, col_reg}<16'b0001011011010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011011010001) && ({row_reg, col_reg}<16'b0001011011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001011011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011011110001) && ({row_reg, col_reg}<16'b0001011011110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011011110100) && ({row_reg, col_reg}<16'b0001011011111011)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0001011011111011) && ({row_reg, col_reg}<16'b0001011100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011100000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001011100000110) && ({row_reg, col_reg}<16'b0001011100001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011100001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011100001011) && ({row_reg, col_reg}<16'b0001011100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011100010010) && ({row_reg, col_reg}<16'b0001011100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001011100100101) && ({row_reg, col_reg}<16'b0001011100100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011100100111) && ({row_reg, col_reg}<16'b0001011100101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011100101011) && ({row_reg, col_reg}<16'b0001011100110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011100110010) && ({row_reg, col_reg}<16'b0001011100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001011100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011100110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001011100111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011100111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001011100111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011100111011) && ({row_reg, col_reg}<16'b0001011101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011101000001) && ({row_reg, col_reg}<16'b0001011101000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001011101000100) && ({row_reg, col_reg}<16'b0001011101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011101000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001011101000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001011101001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001011101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011101001010) && ({row_reg, col_reg}<16'b0001011101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011101001100) && ({row_reg, col_reg}<16'b0001011101010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011101010000) && ({row_reg, col_reg}<16'b0001011101011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011101011000) && ({row_reg, col_reg}<16'b0001011101011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011101011010) && ({row_reg, col_reg}<16'b0001011101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011101011110) && ({row_reg, col_reg}<16'b0001011101100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001011101100001) && ({row_reg, col_reg}<16'b0001011101100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001011101100100) && ({row_reg, col_reg}<16'b0001011101101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001011101101001) && ({row_reg, col_reg}<16'b0001011101101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011101101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001011101101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001011101101101) && ({row_reg, col_reg}<16'b0001011101110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001011101110000) && ({row_reg, col_reg}<16'b0001011101110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001011101110011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0001011101110100) && ({row_reg, col_reg}<16'b0001011101110111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0001011101110111) && ({row_reg, col_reg}<16'b0001011101111100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001011101111100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001011101111101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001011101111110)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0001011101111111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001011110000000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001011110000001) && ({row_reg, col_reg}<16'b0001011110000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011110000011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001011110000100) && ({row_reg, col_reg}<16'b0001011110000110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001011110000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001011110000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011110001000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001011110001001) && ({row_reg, col_reg}<16'b0001011110001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011110001100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001011110001101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001011110001110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001011110001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011110010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011110010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001011110010010) && ({row_reg, col_reg}<16'b0001011110010100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001011110010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001011110010101) && ({row_reg, col_reg}<16'b0001011110011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001011110011000) && ({row_reg, col_reg}<16'b0001011110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001011110011010) && ({row_reg, col_reg}<16'b0001011110011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001011110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001011110011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011110011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011110011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011110100000) && ({row_reg, col_reg}<16'b0001011110100010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001011110100010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0001011110100011) && ({row_reg, col_reg}<16'b0001011110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001011110100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0001011110100111) && ({row_reg, col_reg}<16'b0001011110101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011110101101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001011110101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011110101111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001011110110000) && ({row_reg, col_reg}<16'b0001011110110010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0001011110110010) && ({row_reg, col_reg}<16'b0001011110110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011110110100) && ({row_reg, col_reg}<16'b0001011110110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011110110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001011110111000) && ({row_reg, col_reg}<16'b0001011110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011110111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001011110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001011111000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001011111000001) && ({row_reg, col_reg}<16'b0001011111000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011111000011) && ({row_reg, col_reg}<16'b0001011111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011111000110) && ({row_reg, col_reg}<16'b0001011111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011111001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001011111001001) && ({row_reg, col_reg}<16'b0001011111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011111001011) && ({row_reg, col_reg}<16'b0001011111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011111001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001011111001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011111010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011111010001) && ({row_reg, col_reg}<16'b0001011111101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001011111101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001011111101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001011111101111) && ({row_reg, col_reg}<16'b0001011111110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011111110010) && ({row_reg, col_reg}<16'b0001011111110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011111110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011111111000) && ({row_reg, col_reg}<16'b0001011111111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011111111010)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0001011111111011) && ({row_reg, col_reg}<16'b0001100000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100000000000) && ({row_reg, col_reg}<16'b0001100000000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100000000101) && ({row_reg, col_reg}<16'b0001100000000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100000000111) && ({row_reg, col_reg}<16'b0001100000001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100000001001) && ({row_reg, col_reg}<16'b0001100000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100000010010) && ({row_reg, col_reg}<16'b0001100000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001100000100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100000100110) && ({row_reg, col_reg}<16'b0001100000101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001100000101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001100000101010) && ({row_reg, col_reg}<16'b0001100000101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001100000101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100000101110) && ({row_reg, col_reg}<16'b0001100000110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100000110000) && ({row_reg, col_reg}<16'b0001100000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100000110100) && ({row_reg, col_reg}<16'b0001100000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001100000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100000110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001100000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100000111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001100000111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100000111011) && ({row_reg, col_reg}<16'b0001100001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100001000001) && ({row_reg, col_reg}<16'b0001100001000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001100001000100) && ({row_reg, col_reg}<16'b0001100001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100001000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001100001000111) && ({row_reg, col_reg}<16'b0001100001001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001100001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100001001010) && ({row_reg, col_reg}<16'b0001100001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100001001100) && ({row_reg, col_reg}<16'b0001100001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100001001111) && ({row_reg, col_reg}<16'b0001100001010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100001010111) && ({row_reg, col_reg}<16'b0001100001011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100001011010) && ({row_reg, col_reg}<16'b0001100001011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100001011101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001100001011110) && ({row_reg, col_reg}<16'b0001100001100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100001100001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001100001100010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001100001100011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001100001100100) && ({row_reg, col_reg}<16'b0001100001101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100001101000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001100001101001) && ({row_reg, col_reg}<16'b0001100001101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100001101011) && ({row_reg, col_reg}<16'b0001100001101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100001101101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001100001101110) && ({row_reg, col_reg}<16'b0001100001110000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001100001110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001100001110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100001110010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001100001110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001100001110100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001100001110101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0001100001110110) && ({row_reg, col_reg}<16'b0001100010000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001100010000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001100010000001) && ({row_reg, col_reg}<16'b0001100010000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100010000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100010000100)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0001100010000101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001100010000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001100010000111) && ({row_reg, col_reg}<16'b0001100010001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100010001011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001100010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001100010001101) && ({row_reg, col_reg}<16'b0001100010001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001100010001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001100010010000) && ({row_reg, col_reg}<16'b0001100010010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100010010010) && ({row_reg, col_reg}<16'b0001100010010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001100010010101) && ({row_reg, col_reg}<16'b0001100010011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001100010011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001100010011010) && ({row_reg, col_reg}<16'b0001100010011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001100010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001100010011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100010011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100010011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100010100000) && ({row_reg, col_reg}<16'b0001100010100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001100010100010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0001100010100011) && ({row_reg, col_reg}<16'b0001100010100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001100010100111) && ({row_reg, col_reg}<16'b0001100010110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100010110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001100010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100010110100) && ({row_reg, col_reg}<16'b0001100010110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100010110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001100010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100010111001) && ({row_reg, col_reg}<16'b0001100010111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001100010111011) && ({row_reg, col_reg}<16'b0001100011000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001100011000001) && ({row_reg, col_reg}<16'b0001100011000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100011000011) && ({row_reg, col_reg}<16'b0001100011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100011000110) && ({row_reg, col_reg}<16'b0001100011001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100011001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100011001100) && ({row_reg, col_reg}<16'b0001100011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100011010001) && ({row_reg, col_reg}<16'b0001100011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001100011101101) && ({row_reg, col_reg}<16'b0001100011101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001100011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100011110001) && ({row_reg, col_reg}<16'b0001100011110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100011110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100011111000) && ({row_reg, col_reg}<16'b0001100011111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100011111100) && ({row_reg, col_reg}<16'b0001100011111111)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}==16'b0001100011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001100100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100100000001) && ({row_reg, col_reg}<16'b0001100100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100100000101) && ({row_reg, col_reg}<16'b0001100100000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100100000111) && ({row_reg, col_reg}<16'b0001100100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100100001001) && ({row_reg, col_reg}<16'b0001100100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100100010010) && ({row_reg, col_reg}<16'b0001100100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001100100100101) && ({row_reg, col_reg}<16'b0001100100100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100100100111) && ({row_reg, col_reg}<16'b0001100100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100100101001) && ({row_reg, col_reg}<16'b0001100100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001100100101110) && ({row_reg, col_reg}<16'b0001100100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001100100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100100110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100100110010) && ({row_reg, col_reg}<16'b0001100100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100100110100) && ({row_reg, col_reg}<16'b0001100100110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001100100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100100110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001100100111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100100111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001100100111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001100100111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100100111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001100100111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001100100111110) && ({row_reg, col_reg}<16'b0001100101000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001100101000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100101000001) && ({row_reg, col_reg}<16'b0001100101000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001100101000100) && ({row_reg, col_reg}<16'b0001100101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100101000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001100101000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001100101001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001100101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100101001010) && ({row_reg, col_reg}<16'b0001100101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100101001100) && ({row_reg, col_reg}<16'b0001100101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100101001111) && ({row_reg, col_reg}<16'b0001100101010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100101010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100101010100) && ({row_reg, col_reg}<16'b0001100101010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100101010111) && ({row_reg, col_reg}<16'b0001100101011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100101011010) && ({row_reg, col_reg}<16'b0001100101011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100101011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001100101011110) && ({row_reg, col_reg}<16'b0001100101100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100101100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001100101100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001100101100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001100101100100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001100101100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100101100110) && ({row_reg, col_reg}<16'b0001100101101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001100101101000) && ({row_reg, col_reg}<16'b0001100101101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100101101011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001100101101100) && ({row_reg, col_reg}<16'b0001100101110001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001100101110001) && ({row_reg, col_reg}<16'b0001100101110011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001100101110011) && ({row_reg, col_reg}<16'b0001100101111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001100101111000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0001100101111001) && ({row_reg, col_reg}<16'b0001100101111100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001100101111100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0001100101111101) && ({row_reg, col_reg}<16'b0001100110000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001100110000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100110000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100110000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001100110000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100110000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001100110000101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001100110000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001100110000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100110001000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001100110001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100110001010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001100110001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100110001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100110001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001100110001110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001100110001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100110010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001100110010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001100110010010) && ({row_reg, col_reg}<16'b0001100110010100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001100110010100) && ({row_reg, col_reg}<16'b0001100110010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001100110010110) && ({row_reg, col_reg}<16'b0001100110011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001100110011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001100110011010) && ({row_reg, col_reg}<16'b0001100110011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001100110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001100110011101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001100110011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100110011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100110100000) && ({row_reg, col_reg}<16'b0001100110100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001100110100010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0001100110100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001100110100100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0001100110100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001100110100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100110100111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001100110101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001100110101001) && ({row_reg, col_reg}<16'b0001100110101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100110101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100110101110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001100110101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100110110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001100110110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100110110010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001100110110011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0001100110110100) && ({row_reg, col_reg}<16'b0001100110110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100110110110) && ({row_reg, col_reg}<16'b0001100110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001100110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100110111001) && ({row_reg, col_reg}<16'b0001100110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100110111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001100110111110) && ({row_reg, col_reg}<16'b0001100111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001100111000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001100111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100111000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001100111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001100111000100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100111000101) && ({row_reg, col_reg}<16'b0001100111001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100111001111) && ({row_reg, col_reg}<16'b0001100111010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100111010001) && ({row_reg, col_reg}<16'b0001100111101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001100111101111) && ({row_reg, col_reg}<16'b0001100111110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100111110100) && ({row_reg, col_reg}<16'b0001100111111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100111111000) && ({row_reg, col_reg}<16'b0001100111111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100111111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100111111100) && ({row_reg, col_reg}<16'b0001100111111110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0001100111111110) && ({row_reg, col_reg}<16'b0001101000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101000000001) && ({row_reg, col_reg}<16'b0001101000000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001101000000011) && ({row_reg, col_reg}<16'b0001101000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101000001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101000001110) && ({row_reg, col_reg}<16'b0001101000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101000010010) && ({row_reg, col_reg}<16'b0001101000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001101000100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101000100110) && ({row_reg, col_reg}<16'b0001101000101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101000101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101000101001) && ({row_reg, col_reg}<16'b0001101000101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001101000101110) && ({row_reg, col_reg}<16'b0001101000110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101000110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001101000110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101000110011) && ({row_reg, col_reg}<16'b0001101000110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001101000110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001101000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101000110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001101000111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001101000111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001101000111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101000111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101000111100) && ({row_reg, col_reg}<16'b0001101000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001101000111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101000111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001101001000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001101001000001) && ({row_reg, col_reg}<16'b0001101001000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101001000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001101001000100) && ({row_reg, col_reg}<16'b0001101001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101001000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001101001000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101001001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001101001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001101001001010) && ({row_reg, col_reg}<16'b0001101001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001101001001100) && ({row_reg, col_reg}<16'b0001101001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001101001001110) && ({row_reg, col_reg}<16'b0001101001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101001010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001101001010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101001010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101001010011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0001101001010100) && ({row_reg, col_reg}<16'b0001101001011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001101001011011) && ({row_reg, col_reg}<16'b0001101001011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101001011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001101001011111) && ({row_reg, col_reg}<16'b0001101001100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101001100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001101001100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001101001100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001101001100100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001101001100101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001101001100110) && ({row_reg, col_reg}<16'b0001101001101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101001101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001101001101001) && ({row_reg, col_reg}<16'b0001101001101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101001101011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001101001101100) && ({row_reg, col_reg}<16'b0001101001110001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001101001110001) && ({row_reg, col_reg}<16'b0001101001110011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001101001110011) && ({row_reg, col_reg}<16'b0001101001110111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001101001110111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0001101001111000) && ({row_reg, col_reg}<16'b0001101001111101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001101001111101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001101001111110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001101001111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101010000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101010000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001101010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101010000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101010000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101010000101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0001101010000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001101010000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101010001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101010001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101010001010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001101010001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101010001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001101010001110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001101010001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101010010000)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0001101010010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001101010010010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001101010010011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001101010010100) && ({row_reg, col_reg}<16'b0001101010010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001101010010110) && ({row_reg, col_reg}<16'b0001101010011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001101010011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101010011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101010011010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001101010011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001101010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001101010011101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001101010011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001101010011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101010100000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001101010100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001101010100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101010100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001101010100100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0001101010100101) && ({row_reg, col_reg}<16'b0001101010101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001101010101000) && ({row_reg, col_reg}<16'b0001101010101010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001101010101010) && ({row_reg, col_reg}<16'b0001101010101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001101010101101) && ({row_reg, col_reg}<16'b0001101010101111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001101010101111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001101010110000) && ({row_reg, col_reg}<16'b0001101010110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001101010110010) && ({row_reg, col_reg}<16'b0001101010110100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101010110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101010110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001101010110111) && ({row_reg, col_reg}<16'b0001101010111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101010111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101010111010) && ({row_reg, col_reg}<16'b0001101010111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001101010111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101010111110) && ({row_reg, col_reg}<16'b0001101011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101011000010) && ({row_reg, col_reg}<16'b0001101011000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101011000101) && ({row_reg, col_reg}<16'b0001101011010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101011010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001101011010001) && ({row_reg, col_reg}<16'b0001101011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001101011101111) && ({row_reg, col_reg}<16'b0001101011110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101011110100) && ({row_reg, col_reg}<16'b0001101011111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001101011111000) && ({row_reg, col_reg}<16'b0001101011111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001101011111100) && ({row_reg, col_reg}<16'b0001101011111110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0001101011111110) && ({row_reg, col_reg}<16'b0001101100000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001101100000001) && ({row_reg, col_reg}<16'b0001101100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101100000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001101100000110) && ({row_reg, col_reg}<16'b0001101100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101100010000) && ({row_reg, col_reg}<16'b0001101100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001101100010010) && ({row_reg, col_reg}<16'b0001101100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001101100100101) && ({row_reg, col_reg}<16'b0001101100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101100101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101100101001) && ({row_reg, col_reg}<16'b0001101100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001101100101110) && ({row_reg, col_reg}<16'b0001101100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001101100110000) && ({row_reg, col_reg}<16'b0001101100110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101100110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001101100110011) && ({row_reg, col_reg}<16'b0001101100110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001101100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101100110111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001101100111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001101100111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001101100111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101100111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001101100111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101100111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001101100111110) && ({row_reg, col_reg}<16'b0001101101000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001101101000000) && ({row_reg, col_reg}<16'b0001101101000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001101101000010) && ({row_reg, col_reg}<16'b0001101101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101101000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001101101000111) && ({row_reg, col_reg}<16'b0001101101001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001101101001001) && ({row_reg, col_reg}<16'b0001101101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101101001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101101001101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0001101101001110) && ({row_reg, col_reg}<16'b0001101101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101101010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001101101010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001101101010010) && ({row_reg, col_reg}<16'b0001101101010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001101101010110) && ({row_reg, col_reg}<16'b0001101101011000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001101101011000) && ({row_reg, col_reg}<16'b0001101101011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001101101011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001101101011011) && ({row_reg, col_reg}<16'b0001101101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101101011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001101101011111) && ({row_reg, col_reg}<16'b0001101101100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001101101100001) && ({row_reg, col_reg}<16'b0001101101100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001101101100011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001101101100100) && ({row_reg, col_reg}<16'b0001101101101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101101101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001101101101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101101101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001101101101011) && ({row_reg, col_reg}<16'b0001101101101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001101101101101) && ({row_reg, col_reg}<16'b0001101101110001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001101101110001) && ({row_reg, col_reg}<16'b0001101101110011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001101101110011) && ({row_reg, col_reg}<16'b0001101101110110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001101101110110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0001101101110111) && ({row_reg, col_reg}<16'b0001101101111101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001101101111101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001101101111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101101111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001101110000000) && ({row_reg, col_reg}<16'b0001101110000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001101110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101110000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101110000100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001101110000101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001101110000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001101110000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101110001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001101110001001) && ({row_reg, col_reg}<16'b0001101110001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101110001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101110001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001101110001101) && ({row_reg, col_reg}<16'b0001101110001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001101110001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001101110010000) && ({row_reg, col_reg}<16'b0001101110010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001101110010010) && ({row_reg, col_reg}<16'b0001101110010100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001101110010100) && ({row_reg, col_reg}<16'b0001101110010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001101110010110) && ({row_reg, col_reg}<16'b0001101110011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001101110011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101110011010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001101110011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001101110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001101110011101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001101110011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101110011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001101110100000) && ({row_reg, col_reg}<16'b0001101110100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101110100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001101110100100) && ({row_reg, col_reg}<16'b0001101110101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001101110101000) && ({row_reg, col_reg}<16'b0001101110101010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001101110101010) && ({row_reg, col_reg}<16'b0001101110101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001101110101101) && ({row_reg, col_reg}<16'b0001101110110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101110110000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001101110110001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001101110110010) && ({row_reg, col_reg}<16'b0001101110110100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101110110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101110110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001101110110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001101110111000) && ({row_reg, col_reg}<16'b0001101110111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101110111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101110111011) && ({row_reg, col_reg}<16'b0001101110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001101110111110) && ({row_reg, col_reg}<16'b0001101111000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001101111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101111000001) && ({row_reg, col_reg}<16'b0001101111000100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101111000100) && ({row_reg, col_reg}<16'b0001101111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101111001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101111001111) && ({row_reg, col_reg}<16'b0001101111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101111010001) && ({row_reg, col_reg}<16'b0001101111101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001101111101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101111101111) && ({row_reg, col_reg}<16'b0001101111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101111110010) && ({row_reg, col_reg}<16'b0001101111110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101111110100) && ({row_reg, col_reg}<16'b0001101111110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101111110110) && ({row_reg, col_reg}<16'b0001101111111000)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0001101111111000) && ({row_reg, col_reg}<16'b0001110000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001110000000001) && ({row_reg, col_reg}<16'b0001110000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110000000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001110000000110) && ({row_reg, col_reg}<16'b0001110000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110000001111) && ({row_reg, col_reg}<16'b0001110000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110000010010) && ({row_reg, col_reg}<16'b0001110000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001110000100101) && ({row_reg, col_reg}<16'b0001110000101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110000101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110000101001) && ({row_reg, col_reg}<16'b0001110000101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001110000101110) && ({row_reg, col_reg}<16'b0001110000110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001110000110000) && ({row_reg, col_reg}<16'b0001110000110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110000110011) && ({row_reg, col_reg}<16'b0001110000110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001110000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110000110111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001110000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110000111001) && ({row_reg, col_reg}<16'b0001110000111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001110000111100) && ({row_reg, col_reg}<16'b0001110000111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110000111110) && ({row_reg, col_reg}<16'b0001110001000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110001000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001110001000001) && ({row_reg, col_reg}<16'b0001110001000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110001000100)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}==16'b0001110001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110001000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110001000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110001001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110001001010) && ({row_reg, col_reg}<16'b0001110001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001110001001100) && ({row_reg, col_reg}<16'b0001110001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110001001111) && ({row_reg, col_reg}<16'b0001110001010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001110001010011) && ({row_reg, col_reg}<16'b0001110001010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110001010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110001010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110001010111) && ({row_reg, col_reg}<16'b0001110001011001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001110001011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110001011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110001011011) && ({row_reg, col_reg}<16'b0001110001011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110001011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001110001011111) && ({row_reg, col_reg}<16'b0001110001100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001110001100001) && ({row_reg, col_reg}<16'b0001110001100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001110001100011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001110001100100) && ({row_reg, col_reg}<16'b0001110001100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110001100111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001110001101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001110001101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110001101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110001101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001110001101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110001101101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001110001101110) && ({row_reg, col_reg}<16'b0001110001110001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001110001110001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001110001110010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001110001110011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0001110001110100) && ({row_reg, col_reg}<16'b0001110001110110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001110001110110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0001110001110111) && ({row_reg, col_reg}<16'b0001110001111101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001110001111101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001110001111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110001111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110010000000) && ({row_reg, col_reg}<16'b0001110010000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110010000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110010000100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001110010000101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001110010000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001110010000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110010001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001110010001001) && ({row_reg, col_reg}<16'b0001110010001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110010001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001110010001101) && ({row_reg, col_reg}<16'b0001110010001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001110010001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110010010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001110010010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110010010010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001110010010011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001110010010100) && ({row_reg, col_reg}<16'b0001110010010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001110010010110) && ({row_reg, col_reg}<16'b0001110010011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001110010011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001110010011010) && ({row_reg, col_reg}<16'b0001110010011101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001110010011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001110010011110) && ({row_reg, col_reg}<16'b0001110010100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001110010100000) && ({row_reg, col_reg}<16'b0001110010100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001110010100011) && ({row_reg, col_reg}<16'b0001110010100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001110010100101) && ({row_reg, col_reg}<16'b0001110010101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110010101001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001110010101010) && ({row_reg, col_reg}<16'b0001110010101100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001110010101100) && ({row_reg, col_reg}<16'b0001110010110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110010110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001110010110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110010110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001110010110011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0001110010110100) && ({row_reg, col_reg}<16'b0001110010110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110010110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110010111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110010111001) && ({row_reg, col_reg}<16'b0001110010111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001110010111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001110010111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001110010111110) && ({row_reg, col_reg}<16'b0001110011000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110011000001) && ({row_reg, col_reg}<16'b0001110011000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110011000101) && ({row_reg, col_reg}<16'b0001110011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110011010001) && ({row_reg, col_reg}<16'b0001110011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001110011101110) && ({row_reg, col_reg}<16'b0001110011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001110011110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001110011110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110011110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001110011110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110011110111)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0001110011111000) && ({row_reg, col_reg}<16'b0001110100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001110100000001) && ({row_reg, col_reg}<16'b0001110100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110100000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001110100000110) && ({row_reg, col_reg}<16'b0001110100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110100010010) && ({row_reg, col_reg}<16'b0001110100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001110100100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110100100110) && ({row_reg, col_reg}<16'b0001110100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110100101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110100101001) && ({row_reg, col_reg}<16'b0001110100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001110100101110) && ({row_reg, col_reg}<16'b0001110100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110100110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110100110010) && ({row_reg, col_reg}<16'b0001110100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110100110100) && ({row_reg, col_reg}<16'b0001110100110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001110100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110100110111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001110100111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110100111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110100111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001110100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110100111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110100111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110100111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001110100111111) && ({row_reg, col_reg}<16'b0001110101000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110101000001) && ({row_reg, col_reg}<16'b0001110101000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001110101000011) && ({row_reg, col_reg}<16'b0001110101000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110101000111) && ({row_reg, col_reg}<16'b0001110101001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110101001010) && ({row_reg, col_reg}<16'b0001110101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001110101001100) && ({row_reg, col_reg}<16'b0001110101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110101001111) && ({row_reg, col_reg}<16'b0001110101010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110101010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110101010100) && ({row_reg, col_reg}<16'b0001110101010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001110101010111) && ({row_reg, col_reg}<16'b0001110101011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110101011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110101011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110101011100) && ({row_reg, col_reg}<16'b0001110101011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001110101011111) && ({row_reg, col_reg}<16'b0001110101100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110101100001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001110101100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001110101100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001110101100100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001110101100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110101100110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001110101100111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001110101101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110101101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110101101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110101101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001110101101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110101101101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001110101101110) && ({row_reg, col_reg}<16'b0001110101110010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001110101110010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001110101110011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001110101110100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001110101110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001110101110110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0001110101110111) && ({row_reg, col_reg}<16'b0001110101111101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001110101111101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001110101111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110101111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110110000000) && ({row_reg, col_reg}<16'b0001110110000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110110000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110110000100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001110110000101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001110110000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001110110000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110110001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001110110001001) && ({row_reg, col_reg}<16'b0001110110001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110110001011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001110110001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001110110001101) && ({row_reg, col_reg}<16'b0001110110001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001110110001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110110010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001110110010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001110110010010) && ({row_reg, col_reg}<16'b0001110110010100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001110110010100) && ({row_reg, col_reg}<16'b0001110110010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001110110010110) && ({row_reg, col_reg}<16'b0001110110011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001110110011001) && ({row_reg, col_reg}<16'b0001110110011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110110011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001110110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001110110011101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001110110011110) && ({row_reg, col_reg}<16'b0001110110100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001110110100000) && ({row_reg, col_reg}<16'b0001110110100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110110100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001110110100100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0001110110100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001110110100110) && ({row_reg, col_reg}<16'b0001110110101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110110101001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001110110101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110110101011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001110110101100) && ({row_reg, col_reg}<16'b0001110110101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001110110101111) && ({row_reg, col_reg}<16'b0001110110110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001110110110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001110110110011) && ({row_reg, col_reg}<16'b0001110110110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001110110110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110110110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110110111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110110111001) && ({row_reg, col_reg}<16'b0001110110111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001110110111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001110110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001110110111110) && ({row_reg, col_reg}<16'b0001110111000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110111000001) && ({row_reg, col_reg}<16'b0001110111000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001110111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001110111000100) && ({row_reg, col_reg}<16'b0001110111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001110111000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110111000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001110111001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110111001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001110111001010) && ({row_reg, col_reg}<16'b0001110111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110111010001) && ({row_reg, col_reg}<16'b0001110111101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001110111101110) && ({row_reg, col_reg}<16'b0001110111110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110111110010) && ({row_reg, col_reg}<16'b0001110111110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001110111110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001110111110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001110111110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110111110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001110111111000) && ({row_reg, col_reg}<16'b0001110111111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110111111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001110111111110)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}==16'b0001110111111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001111000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111000000001) && ({row_reg, col_reg}<16'b0001111000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111000000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111000000110) && ({row_reg, col_reg}<16'b0001111000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111000010010) && ({row_reg, col_reg}<16'b0001111000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001111000100101) && ({row_reg, col_reg}<16'b0001111000101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111000101001) && ({row_reg, col_reg}<16'b0001111000101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001111000101110) && ({row_reg, col_reg}<16'b0001111000110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001111000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111000110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001111000110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111000110011) && ({row_reg, col_reg}<16'b0001111000110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001111000110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001111000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111000110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001111000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111000111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001111000111010) && ({row_reg, col_reg}<16'b0001111001000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001111001000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001111001000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001111001000111) && ({row_reg, col_reg}<16'b0001111001001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001111001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001111001001010) && ({row_reg, col_reg}<16'b0001111001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111001001100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0001111001001101) && ({row_reg, col_reg}<16'b0001111001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001111001001111) && ({row_reg, col_reg}<16'b0001111001010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111001010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111001010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001111001010101) && ({row_reg, col_reg}<16'b0001111001010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111001010111) && ({row_reg, col_reg}<16'b0001111001011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001111001011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111001011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001111001011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001111001011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001111001011101) && ({row_reg, col_reg}<16'b0001111001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111001011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111001100000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001111001100001) && ({row_reg, col_reg}<16'b0001111001100011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001111001100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001111001100100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001111001100101) && ({row_reg, col_reg}<16'b0001111001100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111001100111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001111001101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001111001101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111001101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111001101011) && ({row_reg, col_reg}<16'b0001111001101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001111001101101) && ({row_reg, col_reg}<16'b0001111001101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001111001101111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0001111001110000) && ({row_reg, col_reg}<16'b0001111001111011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001111001111011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0001111001111100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001111001111101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0001111001111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111001111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111010000000) && ({row_reg, col_reg}<16'b0001111010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001111010000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111010000100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001111010000101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001111010000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001111010000111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001111010001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111010001001) && ({row_reg, col_reg}<16'b0001111010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111010001100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001111010001101) && ({row_reg, col_reg}<16'b0001111010001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001111010001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001111010010000) && ({row_reg, col_reg}<16'b0001111010010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001111010010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111010010011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001111010010100) && ({row_reg, col_reg}<16'b0001111010010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001111010010110) && ({row_reg, col_reg}<16'b0001111010011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001111010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001111010011011) && ({row_reg, col_reg}<16'b0001111010011101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001111010011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111010011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111010011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111010100000) && ({row_reg, col_reg}<16'b0001111010100010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001111010100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001111010100011) && ({row_reg, col_reg}<16'b0001111010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001111010100110) && ({row_reg, col_reg}<16'b0001111010101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001111010101001) && ({row_reg, col_reg}<16'b0001111010101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001111010101011) && ({row_reg, col_reg}<16'b0001111010110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111010110011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0001111010110100) && ({row_reg, col_reg}<16'b0001111010110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001111010110110) && ({row_reg, col_reg}<16'b0001111010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111010111001) && ({row_reg, col_reg}<16'b0001111010111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001111010111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001111010111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111010111110) && ({row_reg, col_reg}<16'b0001111011000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001111011000000) && ({row_reg, col_reg}<16'b0001111011000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111011000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001111011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001111011000100) && ({row_reg, col_reg}<16'b0001111011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001111011000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111011000111) && ({row_reg, col_reg}<16'b0001111011001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001111011001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001111011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111011001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111011001100) && ({row_reg, col_reg}<16'b0001111011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111011010001) && ({row_reg, col_reg}<16'b0001111011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001111011101111) && ({row_reg, col_reg}<16'b0001111011110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001111011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111011110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111011110011) && ({row_reg, col_reg}<16'b0001111011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001111011110110) && ({row_reg, col_reg}<16'b0001111011111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111011111000) && ({row_reg, col_reg}<16'b0001111011111110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0001111011111110) && ({row_reg, col_reg}<16'b0001111100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111100000000) && ({row_reg, col_reg}<16'b0001111100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111100000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111100000110) && ({row_reg, col_reg}<16'b0001111100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111100010010) && ({row_reg, col_reg}<16'b0001111100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001111100100101) && ({row_reg, col_reg}<16'b0001111100100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111100100111) && ({row_reg, col_reg}<16'b0001111100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111100101001) && ({row_reg, col_reg}<16'b0001111100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001111100101110) && ({row_reg, col_reg}<16'b0001111100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111100110000) && ({row_reg, col_reg}<16'b0001111100110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111100110010) && ({row_reg, col_reg}<16'b0001111100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111100110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001111100110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001111100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111100110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001111100111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001111100111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001111100111010) && ({row_reg, col_reg}<16'b0001111100111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111100111111) && ({row_reg, col_reg}<16'b0001111101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001111101000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001111101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111101000110) && ({row_reg, col_reg}<16'b0001111101001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001111101001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001111101001001) && ({row_reg, col_reg}<16'b0001111101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111101001100) && ({row_reg, col_reg}<16'b0001111101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001111101001111) && ({row_reg, col_reg}<16'b0001111101010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111101010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111101010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001111101010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111101010110) && ({row_reg, col_reg}<16'b0001111101011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001111101011010) && ({row_reg, col_reg}<16'b0001111101011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001111101011100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001111101011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111101011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111101100000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001111101100001) && ({row_reg, col_reg}<16'b0001111101100011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001111101100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001111101100100) && ({row_reg, col_reg}<16'b0001111101100110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001111101100110) && ({row_reg, col_reg}<16'b0001111101101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111101101000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001111101101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111101101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111101101011) && ({row_reg, col_reg}<16'b0001111101101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111101101101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001111101101110) && ({row_reg, col_reg}<16'b0001111101110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001111101110000) && ({row_reg, col_reg}<16'b0001111101110011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0001111101110011) && ({row_reg, col_reg}<16'b0001111101111001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0001111101111001) && ({row_reg, col_reg}<16'b0001111101111011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001111101111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001111101111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111101111101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001111101111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111101111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111110000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111110000001) && ({row_reg, col_reg}<16'b0001111110000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111110000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111110000100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001111110000101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0001111110000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001111110000111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0001111110001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111110001001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001111110001010) && ({row_reg, col_reg}<16'b0001111110001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111110001100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001111110001101) && ({row_reg, col_reg}<16'b0001111110001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001111110001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001111110010000) && ({row_reg, col_reg}<16'b0001111110010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001111110010010) && ({row_reg, col_reg}<16'b0001111110010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001111110010101) && ({row_reg, col_reg}<16'b0001111110011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001111110011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111110011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001111110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111110011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001111110011100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001111110011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111110011110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001111110011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111110100000) && ({row_reg, col_reg}<16'b0001111110100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001111110100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111110100011) && ({row_reg, col_reg}<16'b0001111110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001111110100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111110100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001111110101000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0001111110101001) && ({row_reg, col_reg}<16'b0001111110101100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001111110101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111110101101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001111110101110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001111110101111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001111110110000) && ({row_reg, col_reg}<16'b0001111110110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111110110100) && ({row_reg, col_reg}<16'b0001111110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001111110111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111110111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001111110111011) && ({row_reg, col_reg}<16'b0001111110111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001111110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111110111110) && ({row_reg, col_reg}<16'b0001111111000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001111111000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001111111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111111000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001111111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001111111000100) && ({row_reg, col_reg}<16'b0001111111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001111111000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111111000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001111111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111111001001) && ({row_reg, col_reg}<16'b0001111111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001111111001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001111111001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111111001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001111111001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001111111001111) && ({row_reg, col_reg}<16'b0001111111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111111010001) && ({row_reg, col_reg}<16'b0001111111101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001111111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111111110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001111111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111111110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111111110011) && ({row_reg, col_reg}<16'b0001111111110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001111111110110) && ({row_reg, col_reg}<16'b0001111111111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111111111000) && ({row_reg, col_reg}<16'b0001111111111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111111111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111111111101) && ({row_reg, col_reg}<16'b0001111111111111)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}==16'b0001111111111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010000000000000) && ({row_reg, col_reg}<16'b0010000000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000000000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000000000110) && ({row_reg, col_reg}<16'b0010000000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000000010010) && ({row_reg, col_reg}<16'b0010000000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010000000100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000000100110) && ({row_reg, col_reg}<16'b0010000000101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010000000101001) && ({row_reg, col_reg}<16'b0010000000101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010000000101110) && ({row_reg, col_reg}<16'b0010000000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000000110001) && ({row_reg, col_reg}<16'b0010000000110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010000000110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000000110100) && ({row_reg, col_reg}<16'b0010000000110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010000000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000000110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010000000111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000000111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000000111010) && ({row_reg, col_reg}<16'b0010000000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000000111110) && ({row_reg, col_reg}<16'b0010000001000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000001000010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010000001000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010000001000100) && ({row_reg, col_reg}<16'b0010000001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010000001000111) && ({row_reg, col_reg}<16'b0010000001001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010000001001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000001001010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010000001001011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010000001001100) && ({row_reg, col_reg}<16'b0010000001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010000001001110) && ({row_reg, col_reg}<16'b0010000001010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000001010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000001010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010000001010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000001010110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000001010111) && ({row_reg, col_reg}<16'b0010000001011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010000001011011) && ({row_reg, col_reg}<16'b0010000001011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000001011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000001011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000001011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000001100000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010000001100001) && ({row_reg, col_reg}<16'b0010000001100011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010000001100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010000001100100) && ({row_reg, col_reg}<16'b0010000001100110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010000001100110) && ({row_reg, col_reg}<16'b0010000001101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000001101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000001101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000001101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000001101011) && ({row_reg, col_reg}<16'b0010000001101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000001101101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010000001101110) && ({row_reg, col_reg}<16'b0010000001110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000001110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010000001110001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010000001110010) && ({row_reg, col_reg}<16'b0010000001110100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010000001110100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010000001110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010000001110110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010000001110111) && ({row_reg, col_reg}<16'b0010000001111100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010000001111100) && ({row_reg, col_reg}<16'b0010000001111110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010000001111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000001111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000010000000) && ({row_reg, col_reg}<16'b0010000010000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010000010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000010000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000010000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000010000101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010000010000110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010000010000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000010001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000010001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000010001010) && ({row_reg, col_reg}<16'b0010000010001100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010000010001100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010000010001101) && ({row_reg, col_reg}<16'b0010000010001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010000010001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010000010010000) && ({row_reg, col_reg}<16'b0010000010010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000010010010) && ({row_reg, col_reg}<16'b0010000010010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010000010010100) && ({row_reg, col_reg}<16'b0010000010010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010000010010111) && ({row_reg, col_reg}<16'b0010000010011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000010011001)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010000010011010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010000010011011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0010000010011100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010000010011101)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010000010011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000010011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000010100000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0010000010100001) && ({row_reg, col_reg}<16'b0010000010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000010100011) && ({row_reg, col_reg}<16'b0010000010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010000010100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010000010100111) && ({row_reg, col_reg}<16'b0010000010110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000010110100) && ({row_reg, col_reg}<16'b0010000010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000010111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000010111010) && ({row_reg, col_reg}<16'b0010000010111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000010111100) && ({row_reg, col_reg}<16'b0010000010111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000010111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010000011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000011000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000011000010) && ({row_reg, col_reg}<16'b0010000011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010000011000100) && ({row_reg, col_reg}<16'b0010000011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010000011000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000011000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010000011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000011001001) && ({row_reg, col_reg}<16'b0010000011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010000011001100) && ({row_reg, col_reg}<16'b0010000011001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000011001111) && ({row_reg, col_reg}<16'b0010000011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000011010001) && ({row_reg, col_reg}<16'b0010000011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010000011110000) && ({row_reg, col_reg}<16'b0010000011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000011110010) && ({row_reg, col_reg}<16'b0010000011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010000011110110) && ({row_reg, col_reg}<16'b0010000011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000011111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010000011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010000011111011) && ({row_reg, col_reg}<16'b0010000011111110)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0010000011111110) && ({row_reg, col_reg}<16'b0010000100000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000100000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000100000010) && ({row_reg, col_reg}<16'b0010000100001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000100001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000100001011) && ({row_reg, col_reg}<16'b0010000100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000100010010) && ({row_reg, col_reg}<16'b0010000100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010000100100100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000100100101) && ({row_reg, col_reg}<16'b0010000100100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000100100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000100101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000100101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000100101010) && ({row_reg, col_reg}<16'b0010000100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010000100101110) && ({row_reg, col_reg}<16'b0010000100110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000100110001) && ({row_reg, col_reg}<16'b0010000100110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000100110011) && ({row_reg, col_reg}<16'b0010000100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000100110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010000100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010000100110111) && ({row_reg, col_reg}<16'b0010000100111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000100111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010000100111010) && ({row_reg, col_reg}<16'b0010000100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000100111110) && ({row_reg, col_reg}<16'b0010000101000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010000101000000) && ({row_reg, col_reg}<16'b0010000101000010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010000101000010) && ({row_reg, col_reg}<16'b0010000101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010000101000110) && ({row_reg, col_reg}<16'b0010000101001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000101001001) && ({row_reg, col_reg}<16'b0010000101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000101001100) && ({row_reg, col_reg}<16'b0010000101001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010000101001110) && ({row_reg, col_reg}<16'b0010000101010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000101010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010000101010011) && ({row_reg, col_reg}<16'b0010000101010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010000101010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000101010110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000101010111) && ({row_reg, col_reg}<16'b0010000101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010000101011011) && ({row_reg, col_reg}<16'b0010000101011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000101011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000101011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000101100000)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0010000101100001) && ({row_reg, col_reg}<16'b0010000101100011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0010000101100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010000101100100) && ({row_reg, col_reg}<16'b0010000101100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000101100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010000101101000) && ({row_reg, col_reg}<16'b0010000101101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000101101010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010000101101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010000101101100) && ({row_reg, col_reg}<16'b0010000101110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010000101110001) && ({row_reg, col_reg}<16'b0010000101110011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010000101110011) && ({row_reg, col_reg}<16'b0010000101111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010000101111001) && ({row_reg, col_reg}<16'b0010000101111100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010000101111100) && ({row_reg, col_reg}<16'b0010000101111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000101111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010000110000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000110000001) && ({row_reg, col_reg}<16'b0010000110000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010000110000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000110000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000110000101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010000110000110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010000110000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000110001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000110001001) && ({row_reg, col_reg}<16'b0010000110001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000110001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010000110001101) && ({row_reg, col_reg}<16'b0010000110001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010000110001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010000110010000) && ({row_reg, col_reg}<16'b0010000110010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000110010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010000110010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000110010100) && ({row_reg, col_reg}<16'b0010000110010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010000110010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000110011000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010000110011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010000110011010) && ({row_reg, col_reg}<16'b0010000110011100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010000110011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010000110011101) && ({row_reg, col_reg}<16'b0010000110011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010000110011111) && ({row_reg, col_reg}<16'b0010000110100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000110100011) && ({row_reg, col_reg}<16'b0010000110100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010000110100111) && ({row_reg, col_reg}<16'b0010000110101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000110101100) && ({row_reg, col_reg}<16'b0010000110101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000110101110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0010000110101111) && ({row_reg, col_reg}<16'b0010000110110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000110110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000110110011) && ({row_reg, col_reg}<16'b0010000110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000110111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010000110111001) && ({row_reg, col_reg}<16'b0010000110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000110111110) && ({row_reg, col_reg}<16'b0010000111000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010000111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000111000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000111000010) && ({row_reg, col_reg}<16'b0010000111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010000111000100) && ({row_reg, col_reg}<16'b0010000111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010000111000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000111000111) && ({row_reg, col_reg}<16'b0010000111001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000111001001) && ({row_reg, col_reg}<16'b0010000111001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000111001011) && ({row_reg, col_reg}<16'b0010000111001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010000111001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000111001111) && ({row_reg, col_reg}<16'b0010000111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000111010001) && ({row_reg, col_reg}<16'b0010000111110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010000111110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000111110111) && ({row_reg, col_reg}<16'b0010000111111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000111111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000111111010) && ({row_reg, col_reg}<16'b0010000111111100)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0010000111111100) && ({row_reg, col_reg}<16'b0010001000000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010001000000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001000000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001000000100) && ({row_reg, col_reg}<16'b0010001000000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001000000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001000001000) && ({row_reg, col_reg}<16'b0010001000001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001000001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001000001011) && ({row_reg, col_reg}<16'b0010001000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001000010000) && ({row_reg, col_reg}<16'b0010001000010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001000010010) && ({row_reg, col_reg}<16'b0010001000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010001000100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001000100110) && ({row_reg, col_reg}<16'b0010001000101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001000101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001000101010) && ({row_reg, col_reg}<16'b0010001000101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010001000101110) && ({row_reg, col_reg}<16'b0010001000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001000110001) && ({row_reg, col_reg}<16'b0010001000110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010001000110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001000110100) && ({row_reg, col_reg}<16'b0010001000110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010001000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001000110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001000111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010001000111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001000111011) && ({row_reg, col_reg}<16'b0010001000111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001000111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010001000111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010001000111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010001001000000) && ({row_reg, col_reg}<16'b0010001001000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010001001000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001001000011) && ({row_reg, col_reg}<16'b0010001001000101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010001001000101) && ({row_reg, col_reg}<16'b0010001001001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010001001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010001001001011) && ({row_reg, col_reg}<16'b0010001001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001001001111) && ({row_reg, col_reg}<16'b0010001001010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001001010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001001010011) && ({row_reg, col_reg}<16'b0010001001010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001001010101) && ({row_reg, col_reg}<16'b0010001001010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001001010111) && ({row_reg, col_reg}<16'b0010001001011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010001001011010) && ({row_reg, col_reg}<16'b0010001001011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001001011100) && ({row_reg, col_reg}<16'b0010001001011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001001011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001001011111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010001001100000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001001100001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0010001001100010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001001100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010001001100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001001100101) && ({row_reg, col_reg}<16'b0010001001101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010001001101010) && ({row_reg, col_reg}<16'b0010001001101100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010001001101100) && ({row_reg, col_reg}<16'b0010001001110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001001110000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010001001110001) && ({row_reg, col_reg}<16'b0010001001110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010001001110011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010001001110100) && ({row_reg, col_reg}<16'b0010001001110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001001110111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010001001111000) && ({row_reg, col_reg}<16'b0010001001111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010001001111011) && ({row_reg, col_reg}<16'b0010001010000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001010000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001010000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001010000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010001010000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001010000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001010000101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010001010000110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010001010000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001010001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010001010001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001010001010) && ({row_reg, col_reg}<16'b0010001010001100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010001010001101) && ({row_reg, col_reg}<16'b0010001010001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010001010001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001010010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001010010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010001010010010) && ({row_reg, col_reg}<16'b0010001010010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010001010010100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0010001010010101) && ({row_reg, col_reg}<16'b0010001010010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001010010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001010011000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010001010011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001010011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001010011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010001010011100) && ({row_reg, col_reg}<16'b0010001010011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001010011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010001010011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001010100000) && ({row_reg, col_reg}<16'b0010001010100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001010100010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010001010100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001010100100)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0010001010100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001010100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0010001010100111) && ({row_reg, col_reg}<16'b0010001010101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001010101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001010101101) && ({row_reg, col_reg}<16'b0010001010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001010110100) && ({row_reg, col_reg}<16'b0010001010110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010001010110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001010110111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0010001010111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001010111001) && ({row_reg, col_reg}<16'b0010001010111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001010111110) && ({row_reg, col_reg}<16'b0010001011000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010001011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001011000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001011000010) && ({row_reg, col_reg}<16'b0010001011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010001011000100) && ({row_reg, col_reg}<16'b0010001011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001011001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001011001001) && ({row_reg, col_reg}<16'b0010001011001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010001011001100) && ({row_reg, col_reg}<16'b0010001011001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001011001111) && ({row_reg, col_reg}<16'b0010001011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001011010001) && ({row_reg, col_reg}<16'b0010001011110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010001011110111) && ({row_reg, col_reg}<16'b0010001011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001011111001) && ({row_reg, col_reg}<16'b0010001011111101)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0010001011111101) && ({row_reg, col_reg}<16'b0010001100000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001100000000) && ({row_reg, col_reg}<16'b0010001100000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001100000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001100000100) && ({row_reg, col_reg}<16'b0010001100001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001100001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001100001011) && ({row_reg, col_reg}<16'b0010001100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001100010010) && ({row_reg, col_reg}<16'b0010001100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010001100100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001100100110) && ({row_reg, col_reg}<16'b0010001100101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001100101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001100101011) && ({row_reg, col_reg}<16'b0010001100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010001100101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001100101110) && ({row_reg, col_reg}<16'b0010001100110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001100110001) && ({row_reg, col_reg}<16'b0010001100110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010001100110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001100110100) && ({row_reg, col_reg}<16'b0010001100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001100110110) && ({row_reg, col_reg}<16'b0010001100111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001100111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010001100111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010001100111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001100111100) && ({row_reg, col_reg}<16'b0010001100111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010001100111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010001100111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010001101000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010001101000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001101000010) && ({row_reg, col_reg}<16'b0010001101000101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010001101000101) && ({row_reg, col_reg}<16'b0010001101001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010001101001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010001101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001101001010) && ({row_reg, col_reg}<16'b0010001101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001101001100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0010001101001101) && ({row_reg, col_reg}<16'b0010001101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001101001111) && ({row_reg, col_reg}<16'b0010001101010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001101010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001101010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001101010101) && ({row_reg, col_reg}<16'b0010001101011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001101011000) && ({row_reg, col_reg}<16'b0010001101011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001101011010) && ({row_reg, col_reg}<16'b0010001101011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010001101011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010001101011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001101011110) && ({row_reg, col_reg}<16'b0010001101100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001101100000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001101100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001101100010)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}==16'b0010001101100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001101100100) && ({row_reg, col_reg}<16'b0010001101100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001101100110) && ({row_reg, col_reg}<16'b0010001101101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001101101000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010001101101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001101101010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010001101101011) && ({row_reg, col_reg}<16'b0010001101101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010001101101101) && ({row_reg, col_reg}<16'b0010001101101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001101101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010001101110000) && ({row_reg, col_reg}<16'b0010001101110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010001101110101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010001101110110) && ({row_reg, col_reg}<16'b0010001101111001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010001101111001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0010001101111010) && ({row_reg, col_reg}<16'b0010001101111100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010001101111100) && ({row_reg, col_reg}<16'b0010001101111110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0010001101111110) && ({row_reg, col_reg}<16'b0010001110000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010001110000000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010001110000001) && ({row_reg, col_reg}<16'b0010001110000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001110000100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010001110000101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010001110000110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010001110000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001110001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010001110001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001110001010) && ({row_reg, col_reg}<16'b0010001110001100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001110001100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0010001110001101) && ({row_reg, col_reg}<16'b0010001110001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010001110001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010001110010000) && ({row_reg, col_reg}<16'b0010001110010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010001110010010) && ({row_reg, col_reg}<16'b0010001110010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001110010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010001110010111) && ({row_reg, col_reg}<16'b0010001110011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001110011001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010001110011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001110011011) && ({row_reg, col_reg}<16'b0010001110011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010001110011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001110100000) && ({row_reg, col_reg}<16'b0010001110100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001110100010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010001110100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001110100100)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0010001110100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001110100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0010001110100111) && ({row_reg, col_reg}<16'b0010001110101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010001110101001) && ({row_reg, col_reg}<16'b0010001110101011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010001110101011) && ({row_reg, col_reg}<16'b0010001110101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010001110101101) && ({row_reg, col_reg}<16'b0010001110101111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010001110101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001110110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010001110110001) && ({row_reg, col_reg}<16'b0010001110110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001110110011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010001110110100) && ({row_reg, col_reg}<16'b0010001110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001110111000) && ({row_reg, col_reg}<16'b0010001110111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001110111010) && ({row_reg, col_reg}<16'b0010001110111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010001110111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010001110111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010001111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001111000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001111000010) && ({row_reg, col_reg}<16'b0010001111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010001111000100) && ({row_reg, col_reg}<16'b0010001111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001111000111) && ({row_reg, col_reg}<16'b0010001111001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010001111001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010001111001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001111001011) && ({row_reg, col_reg}<16'b0010001111001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010001111001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010001111001111) && ({row_reg, col_reg}<16'b0010001111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001111010001) && ({row_reg, col_reg}<16'b0010001111110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010001111110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001111111000) && ({row_reg, col_reg}<16'b0010001111111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001111111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010001111111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}==16'b0010001111111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010010000000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010000000001) && ({row_reg, col_reg}<16'b0010010000000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010000000011) && ({row_reg, col_reg}<16'b0010010000000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010000000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010000000110) && ({row_reg, col_reg}<16'b0010010000001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010000001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010010000001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010000001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010000001011) && ({row_reg, col_reg}<16'b0010010000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010000010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010010000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010000010010) && ({row_reg, col_reg}<16'b0010010000100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010010000100110) && ({row_reg, col_reg}<16'b0010010000101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010010000101001) && ({row_reg, col_reg}<16'b0010010000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010000110001) && ({row_reg, col_reg}<16'b0010010000110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010010000110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010000110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010010000110111) && ({row_reg, col_reg}<16'b0010010000111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010000111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010010000111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010000111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010000111100) && ({row_reg, col_reg}<16'b0010010000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010000111110) && ({row_reg, col_reg}<16'b0010010001000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010001000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010001000001) && ({row_reg, col_reg}<16'b0010010001000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010010001000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010001000110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0010010001000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010010001001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010010001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010001001010) && ({row_reg, col_reg}<16'b0010010001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010001001100) && ({row_reg, col_reg}<16'b0010010001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010001001111) && ({row_reg, col_reg}<16'b0010010001010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010001010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010001010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010010001010101) && ({row_reg, col_reg}<16'b0010010001010111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010001010111) && ({row_reg, col_reg}<16'b0010010001011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010001011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010001011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010001011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010010001011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010001011110) && ({row_reg, col_reg}<16'b0010010001100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010001100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010001100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010010001100011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==16'b0010010001100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010001100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010010001100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010001100111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010010001101000) && ({row_reg, col_reg}<16'b0010010001101010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010001101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010010001101011) && ({row_reg, col_reg}<16'b0010010001101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010010001101101) && ({row_reg, col_reg}<16'b0010010001110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010001110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010010001110001) && ({row_reg, col_reg}<16'b0010010001111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010010001111000) && ({row_reg, col_reg}<16'b0010010001111011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010010001111011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0010010001111100) && ({row_reg, col_reg}<16'b0010010001111110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010010001111110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0010010001111111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010010010000000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0010010010000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010010000010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010010010000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010010010000100) && ({row_reg, col_reg}<16'b0010010010000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010010010000110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010010010000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010010001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010010010001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010010001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010010001011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010010010001100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0010010010001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010010010001110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010010010001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010010010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010010010010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010010010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010010010010011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010010010010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010010010101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0010010010010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010010010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010010011000) && ({row_reg, col_reg}<16'b0010010010011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010010011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010010011011) && ({row_reg, col_reg}<16'b0010010010011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010010010011101) && ({row_reg, col_reg}<16'b0010010010011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010010011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010010100000) && ({row_reg, col_reg}<16'b0010010010100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010010100010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010010010100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010010100100)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0010010010100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010010100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0010010010100111) && ({row_reg, col_reg}<16'b0010010010101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010010101011) && ({row_reg, col_reg}<16'b0010010010101101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010010010101101) && ({row_reg, col_reg}<16'b0010010010101111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010010101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010010110000) && ({row_reg, col_reg}<16'b0010010010110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010010110010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010010010110011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010010010110100) && ({row_reg, col_reg}<16'b0010010010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010010111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010010010111011) && ({row_reg, col_reg}<16'b0010010010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010010010111111) && ({row_reg, col_reg}<16'b0010010011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010011000001) && ({row_reg, col_reg}<16'b0010010011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010010011000100) && ({row_reg, col_reg}<16'b0010010011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010011000110) && ({row_reg, col_reg}<16'b0010010011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010011001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010010011001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010010011001010) && ({row_reg, col_reg}<16'b0010010011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010011001111) && ({row_reg, col_reg}<16'b0010010011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010011010001) && ({row_reg, col_reg}<16'b0010010011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010010011110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010011110110) && ({row_reg, col_reg}<16'b0010010011111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010010011111000) && ({row_reg, col_reg}<16'b0010010011111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010011111100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0010010011111101) && ({row_reg, col_reg}<16'b0010010100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010010100000000) && ({row_reg, col_reg}<16'b0010010100000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010010100000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010010100000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010100000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010010100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010100000111) && ({row_reg, col_reg}<16'b0010010100001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010010100001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010100001010) && ({row_reg, col_reg}<16'b0010010100001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010100001100) && ({row_reg, col_reg}<16'b0010010100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010100010010) && ({row_reg, col_reg}<16'b0010010100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010010100100110) && ({row_reg, col_reg}<16'b0010010100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010010100101001) && ({row_reg, col_reg}<16'b0010010100101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010100101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010010100101100) && ({row_reg, col_reg}<16'b0010010100110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010100110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010010100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010010100110011) && ({row_reg, col_reg}<16'b0010010100110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010100110111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010010100111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010010100111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010010100111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010010100111011) && ({row_reg, col_reg}<16'b0010010100111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010100111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010010100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010100111111) && ({row_reg, col_reg}<16'b0010010101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010101000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010010101000010) && ({row_reg, col_reg}<16'b0010010101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010101000100) && ({row_reg, col_reg}<16'b0010010101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010101000111) && ({row_reg, col_reg}<16'b0010010101001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010101001001) && ({row_reg, col_reg}<16'b0010010101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010101001100) && ({row_reg, col_reg}<16'b0010010101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010101001111) && ({row_reg, col_reg}<16'b0010010101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010101010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010101010101) && ({row_reg, col_reg}<16'b0010010101010111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010101010111) && ({row_reg, col_reg}<16'b0010010101011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010101011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010101011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010010101011100) && ({row_reg, col_reg}<16'b0010010101011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010101011110) && ({row_reg, col_reg}<16'b0010010101100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010101100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010101100010) && ({row_reg, col_reg}<16'b0010010101100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010010101100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010101100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010010101100110) && ({row_reg, col_reg}<16'b0010010101101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010101101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010010101101001) && ({row_reg, col_reg}<16'b0010010101101011)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0010010101101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010010101101100) && ({row_reg, col_reg}<16'b0010010101101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010101101111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010010101110000) && ({row_reg, col_reg}<16'b0010010101110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010010101110010) && ({row_reg, col_reg}<16'b0010010101110100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010010101110100) && ({row_reg, col_reg}<16'b0010010101110110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010010101110110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010010101110111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010010101111000) && ({row_reg, col_reg}<16'b0010010101111010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010010101111010)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0010010101111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010010101111100) && ({row_reg, col_reg}<16'b0010010101111110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010010101111110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0010010101111111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010010110000000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0010010110000001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010010110000010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010110000011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010010110000100) && ({row_reg, col_reg}<16'b0010010110000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010010110000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010110000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010110001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010010110001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010110001010) && ({row_reg, col_reg}<16'b0010010110001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010110001100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010010110001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010010110001110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010010110001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010110010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010010110010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010010110010010) && ({row_reg, col_reg}<16'b0010010110010100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010010110010100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010010110010101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0010010110010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010010110010111) && ({row_reg, col_reg}<16'b0010010110011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010110011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010110011011) && ({row_reg, col_reg}<16'b0010010110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010010110011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010110011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010110011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010110100000) && ({row_reg, col_reg}<16'b0010010110100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010110100010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010010110100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010110100100)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}>=16'b0010010110100101) && ({row_reg, col_reg}<16'b0010010110100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010010110100111) && ({row_reg, col_reg}<16'b0010010110101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010110101011) && ({row_reg, col_reg}<16'b0010010110101110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010110101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010010110101111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010010110110000) && ({row_reg, col_reg}<16'b0010010110110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010110110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010110110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010010110111000) && ({row_reg, col_reg}<16'b0010010110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010110111010) && ({row_reg, col_reg}<16'b0010010110111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010010110111100) && ({row_reg, col_reg}<16'b0010010110111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010110111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010010110111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010010111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010111000001) && ({row_reg, col_reg}<16'b0010010111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010010111000100) && ({row_reg, col_reg}<16'b0010010111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010111000110) && ({row_reg, col_reg}<16'b0010010111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010111010001) && ({row_reg, col_reg}<16'b0010010111110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010010111110100) && ({row_reg, col_reg}<16'b0010010111110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010010111110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010111110111) && ({row_reg, col_reg}<16'b0010010111111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010010111111001) && ({row_reg, col_reg}<16'b0010010111111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010111111100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0010010111111101) && ({row_reg, col_reg}<16'b0010011000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011000000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010011000000001) && ({row_reg, col_reg}<16'b0010011000000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011000000011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0010011000000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011000000101) && ({row_reg, col_reg}<16'b0010011000000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010011000000111) && ({row_reg, col_reg}<16'b0010011000001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011000001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010011000001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011000001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011000001101) && ({row_reg, col_reg}<16'b0010011000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011000010010) && ({row_reg, col_reg}<16'b0010011000100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010011000100110) && ({row_reg, col_reg}<16'b0010011000101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010011000101100) && ({row_reg, col_reg}<16'b0010011000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011000110001) && ({row_reg, col_reg}<16'b0010011000110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010011000110100) && ({row_reg, col_reg}<16'b0010011000110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011000110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011000111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010011000111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010011000111010) && ({row_reg, col_reg}<16'b0010011000111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011000111111) && ({row_reg, col_reg}<16'b0010011001000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010011001000010) && ({row_reg, col_reg}<16'b0010011001000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010011001000100) && ({row_reg, col_reg}<16'b0010011001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011001000111) && ({row_reg, col_reg}<16'b0010011001001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010011001001001) && ({row_reg, col_reg}<16'b0010011001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011001001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011001001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011001001110) && ({row_reg, col_reg}<16'b0010011001010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011001010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011001010100) && ({row_reg, col_reg}<16'b0010011001010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011001010110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010011001010111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011001011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011001011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010011001011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010011001011011) && ({row_reg, col_reg}<16'b0010011001011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011001011110) && ({row_reg, col_reg}<16'b0010011001100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011001100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011001100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011001100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010011001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011001100100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010011001100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011001100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011001100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010011001101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011001101001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010011001101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010011001101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010011001101100) && ({row_reg, col_reg}<16'b0010011001101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011001101111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010011001110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010011001110001) && ({row_reg, col_reg}<16'b0010011001110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011001110011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010011001110100) && ({row_reg, col_reg}<16'b0010011001110110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010011001110110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010011001110111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010011001111000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0010011001111001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0010011001111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010011001111011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010011001111100) && ({row_reg, col_reg}<16'b0010011001111110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010011001111110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0010011001111111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010011010000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010011010000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011010000010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010011010000011) && ({row_reg, col_reg}<16'b0010011010000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010011010000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011010000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011010001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011010001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011010001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011010001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011010001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010011010001110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010011010001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011010010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011010010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011010010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010011010010011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010011010010100) && ({row_reg, col_reg}<16'b0010011010010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011010010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010011010010111) && ({row_reg, col_reg}<16'b0010011010011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011010011001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010011010011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011010011011) && ({row_reg, col_reg}<16'b0010011010011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011010011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011010011111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010011010100000) && ({row_reg, col_reg}<16'b0010011010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011010100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011010100100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010011010100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011010101001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010011010101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010011010101011) && ({row_reg, col_reg}<16'b0010011010101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010011010101101) && ({row_reg, col_reg}<16'b0010011010101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011010101111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010011010110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011010110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011010110010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010011010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011010110101) && ({row_reg, col_reg}<16'b0010011010111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010011010111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011010111010) && ({row_reg, col_reg}<16'b0010011010111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010011010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010011010111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011010111110) && ({row_reg, col_reg}<16'b0010011011000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011011000001) && ({row_reg, col_reg}<16'b0010011011000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011011000111) && ({row_reg, col_reg}<16'b0010011011001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011011001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011011001100) && ({row_reg, col_reg}<16'b0010011011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011011010001) && ({row_reg, col_reg}<16'b0010011011110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010011011110100) && ({row_reg, col_reg}<16'b0010011011110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011011110111) && ({row_reg, col_reg}<16'b0010011011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010011011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011011111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011011111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0010011011111100) && ({row_reg, col_reg}<16'b0010011100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010011100000000) && ({row_reg, col_reg}<16'b0010011100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010011100000010) && ({row_reg, col_reg}<16'b0010011100000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011100000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011100001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010011100001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011100001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011100001011) && ({row_reg, col_reg}<16'b0010011100001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011100001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011100001110) && ({row_reg, col_reg}<16'b0010011100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011100010011) && ({row_reg, col_reg}<16'b0010011100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010011100100110) && ({row_reg, col_reg}<16'b0010011100101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010011100101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011100101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011100101110) && ({row_reg, col_reg}<16'b0010011100110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011100110001) && ({row_reg, col_reg}<16'b0010011100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011100110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010011100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011100110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011100111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011100111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010011100111010) && ({row_reg, col_reg}<16'b0010011100111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011100111111) && ({row_reg, col_reg}<16'b0010011101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010011101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011101000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011101001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011101001100) && ({row_reg, col_reg}<16'b0010011101001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010011101001110) && ({row_reg, col_reg}<16'b0010011101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011101010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010011101010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010011101010010) && ({row_reg, col_reg}<16'b0010011101010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011101010100) && ({row_reg, col_reg}<16'b0010011101010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010011101010110) && ({row_reg, col_reg}<16'b0010011101011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011101011000) && ({row_reg, col_reg}<16'b0010011101011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010011101011010) && ({row_reg, col_reg}<16'b0010011101011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011101011111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0010011101100000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011101100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011101100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011101100011) && ({row_reg, col_reg}<16'b0010011101100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011101100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011101100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011101100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011101101000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0010011101101001) && ({row_reg, col_reg}<16'b0010011101101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010011101101011) && ({row_reg, col_reg}<16'b0010011101101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011101101101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0010011101101110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010011101101111) && ({row_reg, col_reg}<16'b0010011101110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011101110011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010011101110100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010011101110101) && ({row_reg, col_reg}<16'b0010011101111000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010011101111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010011101111001) && ({row_reg, col_reg}<16'b0010011101111011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010011101111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010011101111100)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0010011101111101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010011101111110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0010011101111111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010011110000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010011110000001) && ({row_reg, col_reg}<16'b0010011110000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010011110000011) && ({row_reg, col_reg}<16'b0010011110000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010011110000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011110000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011110001000) && ({row_reg, col_reg}<16'b0010011110001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011110001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011110001011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0010011110001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010011110001101) && ({row_reg, col_reg}<16'b0010011110001111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010011110001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010011110010000) && ({row_reg, col_reg}<16'b0010011110010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010011110010010) && ({row_reg, col_reg}<16'b0010011110010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011110010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010011110010101) && ({row_reg, col_reg}<16'b0010011110010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011110010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011110011000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0010011110011001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011110011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011110011011) && ({row_reg, col_reg}<16'b0010011110011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011110011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011110011111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011110100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011110100001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0010011110100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011110100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011110100100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010011110100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010011110100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010011110100111) && ({row_reg, col_reg}<16'b0010011110101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011110101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011110101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010011110101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011110101100) && ({row_reg, col_reg}<16'b0010011110110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010011110110000) && ({row_reg, col_reg}<16'b0010011110110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011110110010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010011110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011110110101) && ({row_reg, col_reg}<16'b0010011110111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010011110111001) && ({row_reg, col_reg}<16'b0010011110111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011110111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010011110111101) && ({row_reg, col_reg}<16'b0010011111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011111000001) && ({row_reg, col_reg}<16'b0010011111000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011111000111) && ({row_reg, col_reg}<16'b0010011111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011111001001) && ({row_reg, col_reg}<16'b0010011111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010011111001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010011111001100) && ({row_reg, col_reg}<16'b0010011111001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010011111001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011111010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011111010001) && ({row_reg, col_reg}<16'b0010011111110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010011111110100) && ({row_reg, col_reg}<16'b0010011111110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011111110111) && ({row_reg, col_reg}<16'b0010011111111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010011111111001) && ({row_reg, col_reg}<16'b0010011111111100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0010011111111100) && ({row_reg, col_reg}<16'b0010100000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100000000001) && ({row_reg, col_reg}<16'b0010100000000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100000000011) && ({row_reg, col_reg}<16'b0010100000000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010100000000111) && ({row_reg, col_reg}<16'b0010100000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010100000001001) && ({row_reg, col_reg}<16'b0010100000001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100000001101) && ({row_reg, col_reg}<16'b0010100000001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100000001111) && ({row_reg, col_reg}<16'b0010100000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100000010010) && ({row_reg, col_reg}<16'b0010100000100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010100000100110) && ({row_reg, col_reg}<16'b0010100000101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100000101100) && ({row_reg, col_reg}<16'b0010100000101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100000101110) && ({row_reg, col_reg}<16'b0010100000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100000110001) && ({row_reg, col_reg}<16'b0010100000110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100000110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010100000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100000110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010100000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100000111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010100000111010) && ({row_reg, col_reg}<16'b0010100000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100000111111) && ({row_reg, col_reg}<16'b0010100001000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100001000100) && ({row_reg, col_reg}<16'b0010100001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100001000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100001000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100001001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010100001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010100001001100) && ({row_reg, col_reg}<16'b0010100001001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010100001001110) && ({row_reg, col_reg}<16'b0010100001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100001010000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010100001010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010100001010010) && ({row_reg, col_reg}<16'b0010100001010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010100001010100) && ({row_reg, col_reg}<16'b0010100001011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010100001011001) && ({row_reg, col_reg}<16'b0010100001011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010100001011011) && ({row_reg, col_reg}<16'b0010100001011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100001011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010100001011111) && ({row_reg, col_reg}<16'b0010100001100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100001100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100001100010) && ({row_reg, col_reg}<16'b0010100001100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100001100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100001100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100001100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010100001101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100001101001)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010100001101010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010100001101011) && ({row_reg, col_reg}<16'b0010100001101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010100001101101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0010100001101110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010100001101111) && ({row_reg, col_reg}<16'b0010100001110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100001110001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010100001110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100001110011) && ({row_reg, col_reg}<16'b0010100001110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010100001110101) && ({row_reg, col_reg}<16'b0010100001111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100001111001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010100001111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100001111011)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0010100001111100) && ({row_reg, col_reg}<16'b0010100001111110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0010100001111110) && ({row_reg, col_reg}<16'b0010100010000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010100010000000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010100010000001) && ({row_reg, col_reg}<16'b0010100010000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100010000011) && ({row_reg, col_reg}<16'b0010100010000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010100010000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100010000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100010001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100010001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010100010001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100010001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100010001100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0010100010001101) && ({row_reg, col_reg}<16'b0010100010001111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010100010001111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010100010010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100010010001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010100010010010) && ({row_reg, col_reg}<16'b0010100010010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100010010100) && ({row_reg, col_reg}<16'b0010100010010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100010010111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010100010011000) && ({row_reg, col_reg}<16'b0010100010011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100010011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100010011011) && ({row_reg, col_reg}<16'b0010100010011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100010011110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010100010011111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010100010100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010100010100001) && ({row_reg, col_reg}<16'b0010100010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100010100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100010100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010100010100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010100010100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010100010101001) && ({row_reg, col_reg}<16'b0010100010101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010100010101100) && ({row_reg, col_reg}<16'b0010100010101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010100010101110) && ({row_reg, col_reg}<16'b0010100010110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100010110100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0010100010110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010100010110110) && ({row_reg, col_reg}<16'b0010100010111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010100010111100) && ({row_reg, col_reg}<16'b0010100010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100010111110) && ({row_reg, col_reg}<16'b0010100011000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100011000001) && ({row_reg, col_reg}<16'b0010100011000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010100011000110) && ({row_reg, col_reg}<16'b0010100011001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100011001011) && ({row_reg, col_reg}<16'b0010100011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010100011001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010100011001111) && ({row_reg, col_reg}<16'b0010100011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100011010001) && ({row_reg, col_reg}<16'b0010100011110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100011110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100011110100) && ({row_reg, col_reg}<16'b0010100011110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100011110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010100011110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100011111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100011111001) && ({row_reg, col_reg}<16'b0010100011111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0010100011111011) && ({row_reg, col_reg}<16'b0010100100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010100100000000) && ({row_reg, col_reg}<16'b0010100100000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010100100000100) && ({row_reg, col_reg}<16'b0010100100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100100000110) && ({row_reg, col_reg}<16'b0010100100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010100100001000) && ({row_reg, col_reg}<16'b0010100100001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010100100001011) && ({row_reg, col_reg}<16'b0010100100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100100001101) && ({row_reg, col_reg}<16'b0010100100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100100010010) && ({row_reg, col_reg}<16'b0010100100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010100100100110) && ({row_reg, col_reg}<16'b0010100100101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100100101100) && ({row_reg, col_reg}<16'b0010100100101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010100100101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100100101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010100100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100100110001) && ({row_reg, col_reg}<16'b0010100100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100100110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010100100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100100110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010100100110111) && ({row_reg, col_reg}<16'b0010100100111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100100111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010100100111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100100111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100100111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100100111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010100100111110) && ({row_reg, col_reg}<16'b0010100101000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100101000000) && ({row_reg, col_reg}<16'b0010100101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010100101000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010100101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100101000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010100101000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010100101001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010100101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010100101001100) && ({row_reg, col_reg}<16'b0010100101001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100101001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010100101001111) && ({row_reg, col_reg}<16'b0010100101010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010100101010011) && ({row_reg, col_reg}<16'b0010100101010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010100101010101) && ({row_reg, col_reg}<16'b0010100101011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010100101011100) && ({row_reg, col_reg}<16'b0010100101011110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010100101011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010100101011111) && ({row_reg, col_reg}<16'b0010100101100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100101100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100101100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100101100011) && ({row_reg, col_reg}<16'b0010100101100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100101100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100101100110) && ({row_reg, col_reg}<16'b0010100101101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100101101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100101101001) && ({row_reg, col_reg}<16'b0010100101101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010100101101101) && ({row_reg, col_reg}<16'b0010100101101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100101101111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010100101110000) && ({row_reg, col_reg}<16'b0010100101110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010100101110011) && ({row_reg, col_reg}<16'b0010100101110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100101110110) && ({row_reg, col_reg}<16'b0010100101111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100101111010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010100101111011) && ({row_reg, col_reg}<16'b0010100110000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100110000011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010100110000100) && ({row_reg, col_reg}<16'b0010100110000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010100110000110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010100110000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100110001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010100110001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100110001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100110001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100110001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100110001101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010100110001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100110001111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010100110010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100110010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100110010010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010100110010011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010100110010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100110010101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010100110010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010100110010111) && ({row_reg, col_reg}<16'b0010100110011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100110011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100110011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100110011100) && ({row_reg, col_reg}<16'b0010100110011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100110011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100110011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010100110100000) && ({row_reg, col_reg}<16'b0010100110100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100110100010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010100110100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100110100100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010100110100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100110100110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010100110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010100110101001) && ({row_reg, col_reg}<16'b0010100110101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100110101011) && ({row_reg, col_reg}<16'b0010100110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100110101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010100110101110) && ({row_reg, col_reg}<16'b0010100110110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010100110110001) && ({row_reg, col_reg}<16'b0010100110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010100110110100) && ({row_reg, col_reg}<16'b0010100110111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100110111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010100110111010) && ({row_reg, col_reg}<16'b0010100110111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100110111100) && ({row_reg, col_reg}<16'b0010100110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100110111110) && ({row_reg, col_reg}<16'b0010100111000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100111000001) && ({row_reg, col_reg}<16'b0010100111000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010100111000110) && ({row_reg, col_reg}<16'b0010100111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100111001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100111001111) && ({row_reg, col_reg}<16'b0010100111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100111010001) && ({row_reg, col_reg}<16'b0010100111110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100111110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100111110101) && ({row_reg, col_reg}<16'b0010100111111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010100111111010)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0010100111111011) && ({row_reg, col_reg}<16'b0010101000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010101000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101000000001) && ({row_reg, col_reg}<16'b0010101000000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010101000000011) && ({row_reg, col_reg}<16'b0010101000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101000000110) && ({row_reg, col_reg}<16'b0010101000001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010101000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010101000001010) && ({row_reg, col_reg}<16'b0010101000010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101000010010) && ({row_reg, col_reg}<16'b0010101000100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010101000100110) && ({row_reg, col_reg}<16'b0010101000101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101000101000) && ({row_reg, col_reg}<16'b0010101000101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101000101011) && ({row_reg, col_reg}<16'b0010101000101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010101000101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101000101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101000110001) && ({row_reg, col_reg}<16'b0010101000110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010101000110100) && ({row_reg, col_reg}<16'b0010101000110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010101000110111) && ({row_reg, col_reg}<16'b0010101000111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101000111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101000111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101000111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010101000111100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101000111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010101000111110) && ({row_reg, col_reg}<16'b0010101001000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101001000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010101001000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101001000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010101001000111) && ({row_reg, col_reg}<16'b0010101001001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010101001001010) && ({row_reg, col_reg}<16'b0010101001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010101001001100) && ({row_reg, col_reg}<16'b0010101001001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010101001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010101001001111) && ({row_reg, col_reg}<16'b0010101001010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101001010010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010101001010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010101001010100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010101001010101) && ({row_reg, col_reg}<16'b0010101001011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101001011001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010101001011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010101001011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101001011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010101001011101)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0010101001011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101001011111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0010101001100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101001100001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010101001100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101001100011) && ({row_reg, col_reg}<16'b0010101001100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010101001100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010101001100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101001100111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010101001101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101001101001)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0010101001101010) && ({row_reg, col_reg}<16'b0010101001101110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010101001101110) && ({row_reg, col_reg}<16'b0010101001110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010101001110000) && ({row_reg, col_reg}<16'b0010101001110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010101001110010) && ({row_reg, col_reg}<16'b0010101001110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010101001110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101001110101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010101001110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101001110111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010101001111000) && ({row_reg, col_reg}<16'b0010101001111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101001111011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0010101001111100) && ({row_reg, col_reg}<16'b0010101001111110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010101001111110) && ({row_reg, col_reg}<16'b0010101010000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101010000001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010101010000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101010000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101010000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101010000101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0010101010000110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010101010000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101010001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101010001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010101010001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010101010001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010101010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101010001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101010001110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010101010001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101010010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010101010010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101010010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101010010011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010101010010100) && ({row_reg, col_reg}<16'b0010101010010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101010010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101010010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010101010011000) && ({row_reg, col_reg}<16'b0010101010011011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010101010011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101010011100) && ({row_reg, col_reg}<16'b0010101010011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010101010011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101010011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101010100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101010100001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010101010100010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010101010100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101010100100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010101010100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101010100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010101010100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010101010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010101010101001) && ({row_reg, col_reg}<16'b0010101010101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101010101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101010101100) && ({row_reg, col_reg}<16'b0010101010101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101010101110) && ({row_reg, col_reg}<16'b0010101010110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010101010110001) && ({row_reg, col_reg}<16'b0010101010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101010110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010101010110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101010110110) && ({row_reg, col_reg}<16'b0010101010111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010101010111000) && ({row_reg, col_reg}<16'b0010101010111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010101010111010) && ({row_reg, col_reg}<16'b0010101010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101010111100) && ({row_reg, col_reg}<16'b0010101010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101010111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010101010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101011000001) && ({row_reg, col_reg}<16'b0010101011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010101011000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101011000110) && ({row_reg, col_reg}<16'b0010101011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101011001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101011001010) && ({row_reg, col_reg}<16'b0010101011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101011010001) && ({row_reg, col_reg}<16'b0010101011110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010101011110100) && ({row_reg, col_reg}<16'b0010101011110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010101011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010101011110111) && ({row_reg, col_reg}<16'b0010101011111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010101011111010)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0010101011111011) && ({row_reg, col_reg}<16'b0010101100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010101100000000) && ({row_reg, col_reg}<16'b0010101100000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010101100000011) && ({row_reg, col_reg}<16'b0010101100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101100000110) && ({row_reg, col_reg}<16'b0010101100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010101100001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101100001001) && ({row_reg, col_reg}<16'b0010101100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101100001101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010101100001110) && ({row_reg, col_reg}<16'b0010101100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101100010010) && ({row_reg, col_reg}<16'b0010101100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010101100100101) && ({row_reg, col_reg}<16'b0010101100101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010101100101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101100101001) && ({row_reg, col_reg}<16'b0010101100101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101100101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101100101100) && ({row_reg, col_reg}<16'b0010101100101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101100101110) && ({row_reg, col_reg}<16'b0010101100110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101100110001) && ({row_reg, col_reg}<16'b0010101100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010101100110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010101100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101100110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010101100110111) && ({row_reg, col_reg}<16'b0010101100111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101100111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101100111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101100111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010101100111100) && ({row_reg, col_reg}<16'b0010101100111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010101100111110) && ({row_reg, col_reg}<16'b0010101101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101101000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010101101000100) && ({row_reg, col_reg}<16'b0010101101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101101000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101101001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010101101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010101101001010) && ({row_reg, col_reg}<16'b0010101101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010101101001100) && ({row_reg, col_reg}<16'b0010101101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010101101001111) && ({row_reg, col_reg}<16'b0010101101010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101101010010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010101101010011)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0010101101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010101101010101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010101101010110) && ({row_reg, col_reg}<16'b0010101101011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101101011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010101101011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010101101011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101101011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010101101011101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010101101011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010101101011111) && ({row_reg, col_reg}<16'b0010101101100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010101101100001) && ({row_reg, col_reg}<16'b0010101101100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101101100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101101100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101101100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010101101100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101101100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101101101000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0010101101101001) && ({row_reg, col_reg}<16'b0010101101101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010101101101011) && ({row_reg, col_reg}<16'b0010101101101110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010101101101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101101101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010101101110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101101110001) && ({row_reg, col_reg}<16'b0010101101110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010101101110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101101110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101101110101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010101101110110) && ({row_reg, col_reg}<16'b0010101101111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101101111100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010101101111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101101111110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010101101111111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101110000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101110000001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010101110000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101110000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010101110000100) && ({row_reg, col_reg}<16'b0010101110000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101110000110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010101110000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101110001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101110001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010101110001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101110001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010101110001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101110001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101110001110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010101110001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101110010000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010101110010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101110010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101110010011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010101110010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101110010101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0010101110010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010101110010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010101110011000) && ({row_reg, col_reg}<16'b0010101110011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010101110011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010101110011011) && ({row_reg, col_reg}<16'b0010101110011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101110011110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010101110011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101110100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101110100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010101110100010) && ({row_reg, col_reg}<16'b0010101110100100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010101110100100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0010101110100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010101110100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010101110100111) && ({row_reg, col_reg}<16'b0010101110101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010101110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101110101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101110101011) && ({row_reg, col_reg}<16'b0010101110101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010101110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101110101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010101110101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010101110110000) && ({row_reg, col_reg}<16'b0010101110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101110110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010101110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101110110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101110110111) && ({row_reg, col_reg}<16'b0010101110111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101110111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010101110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101110111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010101110111100) && ({row_reg, col_reg}<16'b0010101110111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101110111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010101110111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101111000001) && ({row_reg, col_reg}<16'b0010101111000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010101111000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101111000110) && ({row_reg, col_reg}<16'b0010101111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101111010001) && ({row_reg, col_reg}<16'b0010101111110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010101111110100) && ({row_reg, col_reg}<16'b0010101111110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010101111110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101111110111) && ({row_reg, col_reg}<16'b0010101111111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010101111111010)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0010101111111011) && ({row_reg, col_reg}<16'b0010110000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110000000000) && ({row_reg, col_reg}<16'b0010110000000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010110000000010) && ({row_reg, col_reg}<16'b0010110000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110000000110) && ({row_reg, col_reg}<16'b0010110000001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010110000001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110000001001) && ({row_reg, col_reg}<16'b0010110000001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110000001011) && ({row_reg, col_reg}<16'b0010110000001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110000001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010110000001111) && ({row_reg, col_reg}<16'b0010110000010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110000010011) && ({row_reg, col_reg}<16'b0010110000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110000100101) && ({row_reg, col_reg}<16'b0010110000100111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110000100111) && ({row_reg, col_reg}<16'b0010110000101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110000101001) && ({row_reg, col_reg}<16'b0010110000101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110000101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110000101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110000101101) && ({row_reg, col_reg}<16'b0010110000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110000110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110000110001) && ({row_reg, col_reg}<16'b0010110000110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010110000110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010110000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110000110110) && ({row_reg, col_reg}<16'b0010110000111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110000111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110000111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110000111011) && ({row_reg, col_reg}<16'b0010110000111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010110000111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110000111110) && ({row_reg, col_reg}<16'b0010110001000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110001000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110001000100) && ({row_reg, col_reg}<16'b0010110001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110001000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110001001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010110001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010110001001010) && ({row_reg, col_reg}<16'b0010110001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010110001001100) && ({row_reg, col_reg}<16'b0010110001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010110001001110) && ({row_reg, col_reg}<16'b0010110001010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110001010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110001010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010110001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010110001010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010110001010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110001010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010110001011000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010110001011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010110001011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010110001011011) && ({row_reg, col_reg}<16'b0010110001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110001011111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010110001100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110001100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110001100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010110001100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110001100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110001100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110001100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110001100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110001101000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0010110001101001) && ({row_reg, col_reg}<16'b0010110001101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010110001101011) && ({row_reg, col_reg}<16'b0010110001101111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010110001101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110001110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110001110001) && ({row_reg, col_reg}<16'b0010110001110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010110001110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110001110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110001110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010110001110110) && ({row_reg, col_reg}<16'b0010110001111000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010110001111000) && ({row_reg, col_reg}<16'b0010110001111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110001111101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010110001111110) && ({row_reg, col_reg}<16'b0010110010000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010110010000000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010110010000001) && ({row_reg, col_reg}<16'b0010110010000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110010000100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010110010000101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010110010000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110010000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110010001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110010001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010110010001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110010001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010110010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110010001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010110010001110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010110010001111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010110010010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110010010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110010010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010110010010011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010110010010100) && ({row_reg, col_reg}<16'b0010110010010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110010010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010110010010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010110010011000) && ({row_reg, col_reg}<16'b0010110010011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110010011010) && ({row_reg, col_reg}<16'b0010110010011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110010011110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010110010011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010110010100000) && ({row_reg, col_reg}<16'b0010110010100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110010100010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010110010100011) && ({row_reg, col_reg}<16'b0010110010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010110010100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010110010100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110010101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010110010101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110010101010) && ({row_reg, col_reg}<16'b0010110010101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010110010101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110010101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010110010101111) && ({row_reg, col_reg}<16'b0010110010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110010110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110010110101) && ({row_reg, col_reg}<16'b0010110010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110010111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010110010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110010111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110010111100) && ({row_reg, col_reg}<16'b0010110010111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110010111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010110010111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010110011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110011000001) && ({row_reg, col_reg}<16'b0010110011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010110011000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110011000110) && ({row_reg, col_reg}<16'b0010110011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110011001111) && ({row_reg, col_reg}<16'b0010110011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110011010001) && ({row_reg, col_reg}<16'b0010110011110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110011110100) && ({row_reg, col_reg}<16'b0010110011110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010110011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110011110111) && ({row_reg, col_reg}<16'b0010110011111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010110011111010)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0010110011111011) && ({row_reg, col_reg}<16'b0010110100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110100000000) && ({row_reg, col_reg}<16'b0010110100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010110100001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010110100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110100001010) && ({row_reg, col_reg}<16'b0010110100001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110100001110) && ({row_reg, col_reg}<16'b0010110100010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010110100010000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110100010001) && ({row_reg, col_reg}<16'b0010110100010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110100010011) && ({row_reg, col_reg}<16'b0010110100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110100100100) && ({row_reg, col_reg}<16'b0010110100100110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110100100110) && ({row_reg, col_reg}<16'b0010110100101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110100101001) && ({row_reg, col_reg}<16'b0010110100101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110100101011) && ({row_reg, col_reg}<16'b0010110100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110100110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110100110001) && ({row_reg, col_reg}<16'b0010110100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110100110100) && ({row_reg, col_reg}<16'b0010110100110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110100110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110100110111) && ({row_reg, col_reg}<16'b0010110100111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110100111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110100111010) && ({row_reg, col_reg}<16'b0010110100111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110100111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010110100111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110100111110) && ({row_reg, col_reg}<16'b0010110101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110101000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110101000100) && ({row_reg, col_reg}<16'b0010110101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110101000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110101001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010110101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110101001100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010110101001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010110101001110) && ({row_reg, col_reg}<16'b0010110101010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010110101010010) && ({row_reg, col_reg}<16'b0010110101010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010110101010100) && ({row_reg, col_reg}<16'b0010110101010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010110101010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110101010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010110101011000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010110101011001) && ({row_reg, col_reg}<16'b0010110101011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110101011111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010110101100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110101100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110101100010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010110101100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110101100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010110101100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110101100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010110101100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110101101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010110101101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110101101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010110101101100) && ({row_reg, col_reg}<16'b0010110101101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110101101110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010110101101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110101110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010110101110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010110101110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010110101110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010110101110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010110101110101) && ({row_reg, col_reg}<16'b0010110101110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110101110111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010110101111000) && ({row_reg, col_reg}<16'b0010110101111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110101111100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010110101111101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010110101111110)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0010110101111111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010110110000000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010110110000001) && ({row_reg, col_reg}<16'b0010110110000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010110110000100) && ({row_reg, col_reg}<16'b0010110110000110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010110110000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110110000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010110110001000) && ({row_reg, col_reg}<16'b0010110110001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110110001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110110001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110110001101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010110110001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010110110001111) && ({row_reg, col_reg}<16'b0010110110010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110110010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010110110010010) && ({row_reg, col_reg}<16'b0010110110010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110110010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010110110010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110110010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010110110010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110110011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110110011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110110011010) && ({row_reg, col_reg}<16'b0010110110011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110110011110) && ({row_reg, col_reg}<16'b0010110110100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110110100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010110110100100) && ({row_reg, col_reg}<16'b0010110110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010110110100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010110110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110110101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010110110101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110110101010) && ({row_reg, col_reg}<16'b0010110110101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010110110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110110101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110110101111) && ({row_reg, col_reg}<16'b0010110110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110110110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110110110101) && ({row_reg, col_reg}<16'b0010110110110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110110110111) && ({row_reg, col_reg}<16'b0010110110111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010110110111010) && ({row_reg, col_reg}<16'b0010110110111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110110111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010110110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110110111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010110110111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010110111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110111000001) && ({row_reg, col_reg}<16'b0010110111000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010110111000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110111000110) && ({row_reg, col_reg}<16'b0010110111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110111001001) && ({row_reg, col_reg}<16'b0010110111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110111001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110111001100) && ({row_reg, col_reg}<16'b0010110111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110111001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110111001111) && ({row_reg, col_reg}<16'b0010110111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110111010001) && ({row_reg, col_reg}<16'b0010110111110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110111110011) && ({row_reg, col_reg}<16'b0010110111110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010110111110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110111110110) && ({row_reg, col_reg}<16'b0010110111111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110111111000) && ({row_reg, col_reg}<16'b0010110111111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110111111010)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0010110111111011) && ({row_reg, col_reg}<16'b0010111000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010111000000000) && ({row_reg, col_reg}<16'b0010111000000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010111000000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111000000101) && ({row_reg, col_reg}<16'b0010111000001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010111000001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111000001001) && ({row_reg, col_reg}<16'b0010111000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111000001100) && ({row_reg, col_reg}<16'b0010111000001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111000001110) && ({row_reg, col_reg}<16'b0010111000010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111000010000) && ({row_reg, col_reg}<16'b0010111000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111000010011) && ({row_reg, col_reg}<16'b0010111000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010111000100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111000100110) && ({row_reg, col_reg}<16'b0010111000101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111000101001) && ({row_reg, col_reg}<16'b0010111000101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111000101011) && ({row_reg, col_reg}<16'b0010111000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111000110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111000110001) && ({row_reg, col_reg}<16'b0010111000110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010111000110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111000110100) && ({row_reg, col_reg}<16'b0010111000110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010111000110111) && ({row_reg, col_reg}<16'b0010111000111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111000111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111000111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111000111011) && ({row_reg, col_reg}<16'b0010111001000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111001000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010111001000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111001000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010111001000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111001001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010111001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111001001011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0010111001001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010111001001101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010111001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111001001111) && ({row_reg, col_reg}<16'b0010111001010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010111001010011) && ({row_reg, col_reg}<16'b0010111001011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111001011011) && ({row_reg, col_reg}<16'b0010111001011101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010111001011101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010111001011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111001011111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010111001100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111001100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111001100010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010111001100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010111001100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010111001100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111001100110) && ({row_reg, col_reg}<16'b0010111001101001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010111001101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111001101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111001101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010111001101100) && ({row_reg, col_reg}<16'b0010111001101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111001101110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111001101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111001110000) && ({row_reg, col_reg}<16'b0010111001110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111001110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111001110100) && ({row_reg, col_reg}<16'b0010111001110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111001110110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0010111001110111) && ({row_reg, col_reg}<16'b0010111001111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111001111100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010111001111101) && ({row_reg, col_reg}<16'b0010111010000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010111010000000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010111010000001) && ({row_reg, col_reg}<16'b0010111010000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010111010000100) && ({row_reg, col_reg}<16'b0010111010000110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010111010000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111010000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111010001000) && ({row_reg, col_reg}<16'b0010111010001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111010001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010111010001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111010001101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010111010001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010111010001111) && ({row_reg, col_reg}<16'b0010111010010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010111010010101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0010111010010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010111010010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111010011000) && ({row_reg, col_reg}<16'b0010111010011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111010011110) && ({row_reg, col_reg}<16'b0010111010100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010111010100000) && ({row_reg, col_reg}<16'b0010111010100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111010100010) && ({row_reg, col_reg}<16'b0010111010100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010111010100100) && ({row_reg, col_reg}<16'b0010111010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010111010100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010111010100111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0010111010101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111010101001) && ({row_reg, col_reg}<16'b0010111010101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111010101011) && ({row_reg, col_reg}<16'b0010111010101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010111010101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010111010101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111010101111) && ({row_reg, col_reg}<16'b0010111010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111010110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010111010110101) && ({row_reg, col_reg}<16'b0010111010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111010111000) && ({row_reg, col_reg}<16'b0010111010111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010111010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111010111011) && ({row_reg, col_reg}<16'b0010111010111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010111010111111) && ({row_reg, col_reg}<16'b0010111011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111011000001) && ({row_reg, col_reg}<16'b0010111011000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010111011000110) && ({row_reg, col_reg}<16'b0010111011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111011001001) && ({row_reg, col_reg}<16'b0010111011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010111011001100) && ({row_reg, col_reg}<16'b0010111011001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111011001111) && ({row_reg, col_reg}<16'b0010111011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111011010001) && ({row_reg, col_reg}<16'b0010111011110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010111011110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111011110100) && ({row_reg, col_reg}<16'b0010111011110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111011110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111011111000) && ({row_reg, col_reg}<16'b0010111011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111011111011) && ({row_reg, col_reg}<16'b0010111011111111)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}==16'b0010111011111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111100000000) && ({row_reg, col_reg}<16'b0010111100000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010111100000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111100000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010111100000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111100000101) && ({row_reg, col_reg}<16'b0010111100000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010111100000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111100001000) && ({row_reg, col_reg}<16'b0010111100001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010111100001010) && ({row_reg, col_reg}<16'b0010111100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111100001100) && ({row_reg, col_reg}<16'b0010111100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111100001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111100010000) && ({row_reg, col_reg}<16'b0010111100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111100010011) && ({row_reg, col_reg}<16'b0010111100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010111100100101) && ({row_reg, col_reg}<16'b0010111100101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111100101001) && ({row_reg, col_reg}<16'b0010111100101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111100101011) && ({row_reg, col_reg}<16'b0010111100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111100110000) && ({row_reg, col_reg}<16'b0010111100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010111100110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111100110100) && ({row_reg, col_reg}<16'b0010111100110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111100110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010111100110111) && ({row_reg, col_reg}<16'b0010111100111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111100111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111100111010) && ({row_reg, col_reg}<16'b0010111100111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111100111111) && ({row_reg, col_reg}<16'b0010111101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111101000100) && ({row_reg, col_reg}<16'b0010111101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111101000111) && ({row_reg, col_reg}<16'b0010111101001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111101001001) && ({row_reg, col_reg}<16'b0010111101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111101001011) && ({row_reg, col_reg}<16'b0010111101001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111101001110) && ({row_reg, col_reg}<16'b0010111101010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111101010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010111101010011) && ({row_reg, col_reg}<16'b0010111101010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010111101010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111101010110) && ({row_reg, col_reg}<16'b0010111101011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010111101011000) && ({row_reg, col_reg}<16'b0010111101011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010111101011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111101011100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010111101011101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111101011110) && ({row_reg, col_reg}<16'b0010111101100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111101100000) && ({row_reg, col_reg}<16'b0010111101100010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010111101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111101100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010111101100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111101100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111101100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010111101100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111101101000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0010111101101001) && ({row_reg, col_reg}<16'b0010111101101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010111101101011) && ({row_reg, col_reg}<16'b0010111101101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111101101110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111101101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111101110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111101110001) && ({row_reg, col_reg}<16'b0010111101110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111101110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111101110100) && ({row_reg, col_reg}<16'b0010111101110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111101110110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010111101110111) && ({row_reg, col_reg}<16'b0010111101111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111101111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010111101111100) && ({row_reg, col_reg}<16'b0010111110000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010111110000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0010111110000001) && ({row_reg, col_reg}<16'b0010111110000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010111110000100) && ({row_reg, col_reg}<16'b0010111110000110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010111110000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111110000111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010111110001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111110001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111110001010) && ({row_reg, col_reg}<16'b0010111110001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111110001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111110001101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010111110001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111110001111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010111110010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010111110010001) && ({row_reg, col_reg}<16'b0010111110010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111110010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010111110010101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0010111110010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010111110010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111110011000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010111110011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111110011010) && ({row_reg, col_reg}<16'b0010111110011111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010111110011111) && ({row_reg, col_reg}<16'b0010111110100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111110100011) && ({row_reg, col_reg}<16'b0010111110100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010111110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111110101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111110101001) && ({row_reg, col_reg}<16'b0010111110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111110101011) && ({row_reg, col_reg}<16'b0010111110101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010111110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111110101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010111110101111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0010111110110000) && ({row_reg, col_reg}<16'b0010111110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111110110101) && ({row_reg, col_reg}<16'b0010111110111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111110111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010111110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111110111011) && ({row_reg, col_reg}<16'b0010111110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010111110111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111111000001) && ({row_reg, col_reg}<16'b0010111111000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010111111000110) && ({row_reg, col_reg}<16'b0010111111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111111001000) && ({row_reg, col_reg}<16'b0010111111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111111001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010111111001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010111111001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010111111001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010111111001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111111010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111111010001) && ({row_reg, col_reg}<16'b0010111111110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010111111110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111111110100) && ({row_reg, col_reg}<16'b0010111111111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111111111000) && ({row_reg, col_reg}<16'b0010111111111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111111111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111111111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111111111100) && ({row_reg, col_reg}<16'b0010111111111111)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}==16'b0010111111111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011000000000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011000000000001) && ({row_reg, col_reg}<16'b0011000000000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000000000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011000000000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000000000101) && ({row_reg, col_reg}<16'b0011000000001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011000000001000) && ({row_reg, col_reg}<16'b0011000000001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011000000001010) && ({row_reg, col_reg}<16'b0011000000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000000001100) && ({row_reg, col_reg}<16'b0011000000001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000000001110) && ({row_reg, col_reg}<16'b0011000000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011000000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000000010011) && ({row_reg, col_reg}<16'b0011000000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011000000100101) && ({row_reg, col_reg}<16'b0011000000101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000000101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011000000101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000000101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000000101101) && ({row_reg, col_reg}<16'b0011000000101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000000101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000000110000) && ({row_reg, col_reg}<16'b0011000000110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011000000110010) && ({row_reg, col_reg}<16'b0011000000110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000000110100) && ({row_reg, col_reg}<16'b0011000000110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011000000110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011000000111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011000000111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000000111010) && ({row_reg, col_reg}<16'b0011000000111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000000111111) && ({row_reg, col_reg}<16'b0011000001000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011000001000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011000001000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000001000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011000001000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000001001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011000001001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011000001001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000001001011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0011000001001100) && ({row_reg, col_reg}<16'b0011000001001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011000001001111) && ({row_reg, col_reg}<16'b0011000001010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011000001010001) && ({row_reg, col_reg}<16'b0011000001010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011000001010011) && ({row_reg, col_reg}<16'b0011000001010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011000001010101) && ({row_reg, col_reg}<16'b0011000001011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011000001011000) && ({row_reg, col_reg}<16'b0011000001011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011000001011010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011000001011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011000001011100) && ({row_reg, col_reg}<16'b0011000001011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011000001011110) && ({row_reg, col_reg}<16'b0011000001100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000001100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000001100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011000001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011000001100011) && ({row_reg, col_reg}<16'b0011000001100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000001100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000001100110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011000001100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011000001101000) && ({row_reg, col_reg}<16'b0011000001101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000001101010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011000001101011) && ({row_reg, col_reg}<16'b0011000001101101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011000001101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000001101110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011000001101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000001110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011000001110001) && ({row_reg, col_reg}<16'b0011000001110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011000001110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011000001110100) && ({row_reg, col_reg}<16'b0011000001110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000001110110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0011000001110111) && ({row_reg, col_reg}<16'b0011000001111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000001111011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0011000001111100) && ({row_reg, col_reg}<16'b0011000001111111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011000001111111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011000010000000)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0011000010000001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011000010000010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011000010000011) && ({row_reg, col_reg}<16'b0011000010000110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011000010000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000010000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000010001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000010001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011000010001010) && ({row_reg, col_reg}<16'b0011000010001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000010001101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011000010001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000010001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000010010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000010010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011000010010010) && ({row_reg, col_reg}<16'b0011000010010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011000010010100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0011000010010101) && ({row_reg, col_reg}<16'b0011000010010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011000010010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000010011000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0011000010011001) && ({row_reg, col_reg}<16'b0011000010011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000010011110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011000010011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000010100000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0011000010100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011000010100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011000010100011) && ({row_reg, col_reg}<16'b0011000010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011000010100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000010101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011000010101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000010101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000010101011) && ({row_reg, col_reg}<16'b0011000010101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011000010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000010101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011000010101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011000010110000) && ({row_reg, col_reg}<16'b0011000010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000010110101)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b0011000010110110) && ({row_reg, col_reg}<16'b0011000010111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011000010111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011000010111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011000010111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000010111100) && ({row_reg, col_reg}<16'b0011000010111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011000010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000010111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011000011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000011000001) && ({row_reg, col_reg}<16'b0011000011000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011000011000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000011000111) && ({row_reg, col_reg}<16'b0011000011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000011001011) && ({row_reg, col_reg}<16'b0011000011001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011000011001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000011010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000011010001) && ({row_reg, col_reg}<16'b0011000011110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011000011110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000011110100) && ({row_reg, col_reg}<16'b0011000011110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000011110111) && ({row_reg, col_reg}<16'b0011000011111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011000011111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000011111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000011111100) && ({row_reg, col_reg}<16'b0011000011111111)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}==16'b0011000011111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011000100000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011000100000001) && ({row_reg, col_reg}<16'b0011000100000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000100000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011000100000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000100000101) && ({row_reg, col_reg}<16'b0011000100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011000100001000) && ({row_reg, col_reg}<16'b0011000100001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011000100001010) && ({row_reg, col_reg}<16'b0011000100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000100001100) && ({row_reg, col_reg}<16'b0011000100001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000100001110) && ({row_reg, col_reg}<16'b0011000100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011000100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000100010011) && ({row_reg, col_reg}<16'b0011000100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011000100100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000100100110) && ({row_reg, col_reg}<16'b0011000100101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000100101100) && ({row_reg, col_reg}<16'b0011000100101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011000100101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000100101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000100110000) && ({row_reg, col_reg}<16'b0011000100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011000100110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000100110011) && ({row_reg, col_reg}<16'b0011000100110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000100110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011000100110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011000100111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011000100111001) && ({row_reg, col_reg}<16'b0011000100111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000100111100) && ({row_reg, col_reg}<16'b0011000100111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011000100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000100111111) && ({row_reg, col_reg}<16'b0011000101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011000101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011000101000111) && ({row_reg, col_reg}<16'b0011000101001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000101001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011000101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011000101001100) && ({row_reg, col_reg}<16'b0011000101001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011000101001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011000101001111) && ({row_reg, col_reg}<16'b0011000101010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000101010010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011000101010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011000101010100) && ({row_reg, col_reg}<16'b0011000101011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011000101011000) && ({row_reg, col_reg}<16'b0011000101011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011000101011010) && ({row_reg, col_reg}<16'b0011000101011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000101011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000101011101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011000101011110) && ({row_reg, col_reg}<16'b0011000101100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011000101100001) && ({row_reg, col_reg}<16'b0011000101100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011000101100011) && ({row_reg, col_reg}<16'b0011000101100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011000101100110) && ({row_reg, col_reg}<16'b0011000101101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000101101000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011000101101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000101101010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011000101101011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011000101101100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0011000101101101) && ({row_reg, col_reg}<16'b0011000101101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000101101111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011000101110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011000101110001) && ({row_reg, col_reg}<16'b0011000101110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000101110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000101110101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011000101110110) && ({row_reg, col_reg}<16'b0011000101111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000101111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0011000101111100) && ({row_reg, col_reg}<16'b0011000101111111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011000101111111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011000110000000) && ({row_reg, col_reg}<16'b0011000110000010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011000110000010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000110000011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011000110000100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011000110000101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011000110000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000110000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000110001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011000110001001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0011000110001010) && ({row_reg, col_reg}<16'b0011000110001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000110001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000110001101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011000110001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000110001111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0011000110010000) && ({row_reg, col_reg}<16'b0011000110010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011000110010010) && ({row_reg, col_reg}<16'b0011000110010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000110010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011000110010110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0011000110010111) && ({row_reg, col_reg}<16'b0011000110011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000110011010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011000110011011) && ({row_reg, col_reg}<16'b0011000110011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011000110011101) && ({row_reg, col_reg}<16'b0011000110100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000110100001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0011000110100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000110100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011000110100100) && ({row_reg, col_reg}<16'b0011000110100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011000110101001) && ({row_reg, col_reg}<16'b0011000110101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011000110101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000110101100) && ({row_reg, col_reg}<16'b0011000110101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000110101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011000110101111) && ({row_reg, col_reg}<16'b0011000110110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011000110110001) && ({row_reg, col_reg}<16'b0011000110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000110110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011000110110101)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}>=16'b0011000110110110) && ({row_reg, col_reg}<16'b0011000110111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011000110111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000110111101) && ({row_reg, col_reg}<16'b0011000111000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011000111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000111000001) && ({row_reg, col_reg}<16'b0011000111000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011000111000110) && ({row_reg, col_reg}<16'b0011000111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000111001001) && ({row_reg, col_reg}<16'b0011000111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000111001011) && ({row_reg, col_reg}<16'b0011000111001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000111001111) && ({row_reg, col_reg}<16'b0011000111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000111010001) && ({row_reg, col_reg}<16'b0011000111110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011000111110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000111110100) && ({row_reg, col_reg}<16'b0011000111111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000111111000) && ({row_reg, col_reg}<16'b0011000111111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000111111011) && ({row_reg, col_reg}<16'b0011000111111111)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}==16'b0011000111111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001000000000) && ({row_reg, col_reg}<16'b0011001000000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011001000000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011001000000100) && ({row_reg, col_reg}<16'b0011001000001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001000001000) && ({row_reg, col_reg}<16'b0011001000001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011001000001010) && ({row_reg, col_reg}<16'b0011001000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001000001100) && ({row_reg, col_reg}<16'b0011001000001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001000001110) && ({row_reg, col_reg}<16'b0011001000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011001000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001000010011) && ({row_reg, col_reg}<16'b0011001000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011001000100101) && ({row_reg, col_reg}<16'b0011001000101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011001000101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001000101001) && ({row_reg, col_reg}<16'b0011001000101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011001000101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001000101100) && ({row_reg, col_reg}<16'b0011001000101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001000101110) && ({row_reg, col_reg}<16'b0011001000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001000110000) && ({row_reg, col_reg}<16'b0011001000110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011001000110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011001000110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001000110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011001000110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011001000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011001000110111) && ({row_reg, col_reg}<16'b0011001000111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011001000111001) && ({row_reg, col_reg}<16'b0011001000111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001000111011) && ({row_reg, col_reg}<16'b0011001000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011001000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001000111111) && ({row_reg, col_reg}<16'b0011001001000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011001001000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011001001000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011001001000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011001001000111) && ({row_reg, col_reg}<16'b0011001001001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001001001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011001001001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011001001001011) && ({row_reg, col_reg}<16'b0011001001001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011001001001101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011001001001110) && ({row_reg, col_reg}<16'b0011001001010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001001010010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011001001010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011001001010100) && ({row_reg, col_reg}<16'b0011001001010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001001010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011001001010111) && ({row_reg, col_reg}<16'b0011001001011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001001011001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011001001011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001001011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011001001011100) && ({row_reg, col_reg}<16'b0011001001011110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011001001011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001001011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011001001100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011001001100001) && ({row_reg, col_reg}<16'b0011001001100011)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0011001001100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011001001100100) && ({row_reg, col_reg}<16'b0011001001100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001001100110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011001001100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001001101000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011001001101001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011001001101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011001001101011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011001001101100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011001001101101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011001001101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001001101111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011001001110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001001110001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011001001110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011001001110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011001001110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001001110101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0011001001110110) && ({row_reg, col_reg}<16'b0011001001111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011001001111111) && ({row_reg, col_reg}<16'b0011001010000001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011001010000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011001010000010) && ({row_reg, col_reg}<16'b0011001010000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001010000100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0011001010000101) && ({row_reg, col_reg}<16'b0011001010000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001010000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001010001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011001010001001) && ({row_reg, col_reg}<16'b0011001010001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001010001101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011001010001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011001010001111) && ({row_reg, col_reg}<16'b0011001010010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011001010010010) && ({row_reg, col_reg}<16'b0011001010010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011001010010101) && ({row_reg, col_reg}<16'b0011001010010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011001010010111) && ({row_reg, col_reg}<16'b0011001010011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011001010011010) && ({row_reg, col_reg}<16'b0011001010011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011001010011100) && ({row_reg, col_reg}<16'b0011001010100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001010100001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0011001010100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011001010100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011001010100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001010100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011001010100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011001010101001) && ({row_reg, col_reg}<16'b0011001010101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001010101011) && ({row_reg, col_reg}<16'b0011001010101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001010101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011001010101111) && ({row_reg, col_reg}<16'b0011001010110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011001010110001) && ({row_reg, col_reg}<16'b0011001010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011001010110101) && ({row_reg, col_reg}<16'b0011001010111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001010111011) && ({row_reg, col_reg}<16'b0011001010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001010111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011001010111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011001011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001011000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001011000010) && ({row_reg, col_reg}<16'b0011001011000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011001011000110) && ({row_reg, col_reg}<16'b0011001011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001011001001) && ({row_reg, col_reg}<16'b0011001011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001011001011) && ({row_reg, col_reg}<16'b0011001011001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001011001111) && ({row_reg, col_reg}<16'b0011001011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001011010001) && ({row_reg, col_reg}<16'b0011001011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011001011110000) && ({row_reg, col_reg}<16'b0011001011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001011110010) && ({row_reg, col_reg}<16'b0011001011110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001011110100) && ({row_reg, col_reg}<16'b0011001011110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001011110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001011110111) && ({row_reg, col_reg}<16'b0011001011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011001011111001) && ({row_reg, col_reg}<16'b0011001011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001011111011) && ({row_reg, col_reg}<16'b0011001011111111)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}==16'b0011001011111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001100000000) && ({row_reg, col_reg}<16'b0011001100000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011001100000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011001100000100) && ({row_reg, col_reg}<16'b0011001100001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001100001000) && ({row_reg, col_reg}<16'b0011001100001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011001100001010) && ({row_reg, col_reg}<16'b0011001100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001100001100) && ({row_reg, col_reg}<16'b0011001100001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001100001110) && ({row_reg, col_reg}<16'b0011001100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011001100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001100010011) && ({row_reg, col_reg}<16'b0011001100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011001100100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001100100110) && ({row_reg, col_reg}<16'b0011001100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001100101000) && ({row_reg, col_reg}<16'b0011001100101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001100101110) && ({row_reg, col_reg}<16'b0011001100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001100110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011001100110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011001100110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011001100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001100110100) && ({row_reg, col_reg}<16'b0011001100110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011001100110110) && ({row_reg, col_reg}<16'b0011001100111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011001100111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011001100111001) && ({row_reg, col_reg}<16'b0011001100111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001100111100) && ({row_reg, col_reg}<16'b0011001100111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011001100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001100111111) && ({row_reg, col_reg}<16'b0011001101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001101000100) && ({row_reg, col_reg}<16'b0011001101000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011001101000111) && ({row_reg, col_reg}<16'b0011001101001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001101001001) && ({row_reg, col_reg}<16'b0011001101001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001101001011) && ({row_reg, col_reg}<16'b0011001101001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001101001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011001101001110) && ({row_reg, col_reg}<16'b0011001101010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001101010010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011001101010011) && ({row_reg, col_reg}<16'b0011001101010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011001101010110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011001101010111) && ({row_reg, col_reg}<16'b0011001101011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001101011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011001101011011) && ({row_reg, col_reg}<16'b0011001101011110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011001101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011001101011111) && ({row_reg, col_reg}<16'b0011001101100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011001101100001) && ({row_reg, col_reg}<16'b0011001101100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011001101100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001101100100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011001101100101) && ({row_reg, col_reg}<16'b0011001101100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001101100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011001101101000) && ({row_reg, col_reg}<16'b0011001101101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001101101010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011001101101011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011001101101100)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0011001101101101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011001101101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001101101111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011001101110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001101110001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011001101110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011001101110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011001101110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011001101110101) && ({row_reg, col_reg}<16'b0011001101111000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011001101111000) && ({row_reg, col_reg}<16'b0011001101111010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0011001101111010) && ({row_reg, col_reg}<16'b0011001101111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011001101111100) && ({row_reg, col_reg}<16'b0011001101111111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011001101111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011001110000000) && ({row_reg, col_reg}<16'b0011001110000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001110000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011001110000011) && ({row_reg, col_reg}<16'b0011001110000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011001110000111) && ({row_reg, col_reg}<16'b0011001110001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011001110001001) && ({row_reg, col_reg}<16'b0011001110001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001110001110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011001110001111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011001110010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001110010001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011001110010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001110010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011001110010100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0011001110010101) && ({row_reg, col_reg}<16'b0011001110010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011001110010111) && ({row_reg, col_reg}<16'b0011001110011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011001110011010) && ({row_reg, col_reg}<16'b0011001110011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011001110011101) && ({row_reg, col_reg}<16'b0011001110100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001110100001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0011001110100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011001110100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011001110100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001110100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011001110100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011001110101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011001110101010) && ({row_reg, col_reg}<16'b0011001110101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001110101100) && ({row_reg, col_reg}<16'b0011001110101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011001110101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011001110101111) && ({row_reg, col_reg}<16'b0011001110110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011001110110001) && ({row_reg, col_reg}<16'b0011001110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011001110110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011001110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011001110110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011001110110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011001110111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011001110111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001110111010) && ({row_reg, col_reg}<16'b0011001110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001110111110) && ({row_reg, col_reg}<16'b0011001111000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011001111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001111000001) && ({row_reg, col_reg}<16'b0011001111000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001111000011) && ({row_reg, col_reg}<16'b0011001111000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011001111000101) && ({row_reg, col_reg}<16'b0011001111000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001111000111) && ({row_reg, col_reg}<16'b0011001111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001111001001) && ({row_reg, col_reg}<16'b0011001111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001111001011) && ({row_reg, col_reg}<16'b0011001111001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001111001101) && ({row_reg, col_reg}<16'b0011001111001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011001111001111) && ({row_reg, col_reg}<16'b0011001111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001111010001) && ({row_reg, col_reg}<16'b0011001111101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011001111101111) && ({row_reg, col_reg}<16'b0011001111110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001111110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001111110110) && ({row_reg, col_reg}<16'b0011001111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011001111111001) && ({row_reg, col_reg}<16'b0011001111111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001111111011) && ({row_reg, col_reg}<16'b0011001111111111)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}==16'b0011001111111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010000000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011010000000001) && ({row_reg, col_reg}<16'b0011010000000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010000000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011010000000100) && ({row_reg, col_reg}<16'b0011010000001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010000001000) && ({row_reg, col_reg}<16'b0011010000001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011010000001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011010000001100) && ({row_reg, col_reg}<16'b0011010000001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010000001110) && ({row_reg, col_reg}<16'b0011010000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010000010011) && ({row_reg, col_reg}<16'b0011010000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011010000100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010000100110) && ({row_reg, col_reg}<16'b0011010000101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010000101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010000101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011010000101010) && ({row_reg, col_reg}<16'b0011010000101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010000101110) && ({row_reg, col_reg}<16'b0011010000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010000110000) && ({row_reg, col_reg}<16'b0011010000110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010000110010) && ({row_reg, col_reg}<16'b0011010000110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010000110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010000110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011010000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010000110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011010000111001) && ({row_reg, col_reg}<16'b0011010000111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010000111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011010000111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011010000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010000111111) && ({row_reg, col_reg}<16'b0011010001000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010001000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011010001000100) && ({row_reg, col_reg}<16'b0011010001000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011010001000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010001000111) && ({row_reg, col_reg}<16'b0011010001001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011010001001001) && ({row_reg, col_reg}<16'b0011010001001100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011010001001100) && ({row_reg, col_reg}<16'b0011010001001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011010001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011010001001111) && ({row_reg, col_reg}<16'b0011010001010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010001010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011010001010011) && ({row_reg, col_reg}<16'b0011010001010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011010001010101) && ({row_reg, col_reg}<16'b0011010001010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011010001010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011010001011000) && ({row_reg, col_reg}<16'b0011010001011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010001011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011010001011011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011010001011100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011010001011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010001011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010001011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010001100000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011010001100001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0011010001100010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0011010001100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011010001100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011010001100101) && ({row_reg, col_reg}<16'b0011010001100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010001100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010001101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010001101001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011010001101010)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0011010001101011) && ({row_reg, col_reg}<16'b0011010001101110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011010001101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010001101111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011010001110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011010001110001) && ({row_reg, col_reg}<16'b0011010001110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011010001110011) && ({row_reg, col_reg}<16'b0011010001110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011010001110101) && ({row_reg, col_reg}<16'b0011010001110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010001110111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0011010001111000) && ({row_reg, col_reg}<16'b0011010001111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011010001111010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0011010001111011) && ({row_reg, col_reg}<16'b0011010001111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010001111101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011010001111110)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0011010001111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010010000000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011010010000001) && ({row_reg, col_reg}<16'b0011010010000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011010010000011) && ({row_reg, col_reg}<16'b0011010010000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010010000101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011010010000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010010000111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011010010001000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011010010001001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011010010001010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0011010010001011) && ({row_reg, col_reg}<16'b0011010010001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010010001110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011010010001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011010010010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010010010001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0011010010010010) && ({row_reg, col_reg}<16'b0011010010010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011010010010101) && ({row_reg, col_reg}<16'b0011010010010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011010010010111) && ({row_reg, col_reg}<16'b0011010010011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011010010011011) && ({row_reg, col_reg}<16'b0011010010011101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011010010011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011010010011110) && ({row_reg, col_reg}<16'b0011010010100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010010100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010010100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011010010100100) && ({row_reg, col_reg}<16'b0011010010100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010010101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011010010101010) && ({row_reg, col_reg}<16'b0011010010101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010010101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010010101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011010010101110) && ({row_reg, col_reg}<16'b0011010010110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011010010110000) && ({row_reg, col_reg}<16'b0011010010110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011010010110100) && ({row_reg, col_reg}<16'b0011010010110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011010010110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011010010110111) && ({row_reg, col_reg}<16'b0011010010111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011010010111001) && ({row_reg, col_reg}<16'b0011010010111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011010010111011) && ({row_reg, col_reg}<16'b0011010010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010010111110) && ({row_reg, col_reg}<16'b0011010011000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011010011000000) && ({row_reg, col_reg}<16'b0011010011000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010011000100) && ({row_reg, col_reg}<16'b0011010011001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010011001000) && ({row_reg, col_reg}<16'b0011010011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010011001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010011001100) && ({row_reg, col_reg}<16'b0011010011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010011010001) && ({row_reg, col_reg}<16'b0011010011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011010011101111) && ({row_reg, col_reg}<16'b0011010011110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010011110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010011110110) && ({row_reg, col_reg}<16'b0011010011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011010011111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011010011111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010011111011) && ({row_reg, col_reg}<16'b0011010011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011010011111110)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}==16'b0011010011111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010100000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011010100000001) && ({row_reg, col_reg}<16'b0011010100000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010100000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011010100000100) && ({row_reg, col_reg}<16'b0011010100001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010100001000) && ({row_reg, col_reg}<16'b0011010100001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011010100001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010100001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011010100001100) && ({row_reg, col_reg}<16'b0011010100001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010100001110) && ({row_reg, col_reg}<16'b0011010100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010100010011) && ({row_reg, col_reg}<16'b0011010100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011010100100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010100100110) && ({row_reg, col_reg}<16'b0011010100101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010100101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010100101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011010100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011010100101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010100101110) && ({row_reg, col_reg}<16'b0011010100110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010100110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010100110010) && ({row_reg, col_reg}<16'b0011010100110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010100110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011010100110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011010100110110) && ({row_reg, col_reg}<16'b0011010100111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011010100111001) && ({row_reg, col_reg}<16'b0011010100111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011010100111100) && ({row_reg, col_reg}<16'b0011010100111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011010100111110) && ({row_reg, col_reg}<16'b0011010101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011010101000011) && ({row_reg, col_reg}<16'b0011010101000101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011010101000101) && ({row_reg, col_reg}<16'b0011010101000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011010101000111) && ({row_reg, col_reg}<16'b0011010101001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011010101001100) && ({row_reg, col_reg}<16'b0011010101001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011010101001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011010101001111) && ({row_reg, col_reg}<16'b0011010101010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011010101010010) && ({row_reg, col_reg}<16'b0011010101010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010101010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010101010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011010101010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011010101011000) && ({row_reg, col_reg}<16'b0011010101011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010101011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011010101100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010101100001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0011010101100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011010101100011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0011010101100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011010101100101) && ({row_reg, col_reg}<16'b0011010101100111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011010101100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010101101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011010101101001)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0011010101101010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011010101101011) && ({row_reg, col_reg}<16'b0011010101101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010101101101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011010101101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010101101111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011010101110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011010101110001) && ({row_reg, col_reg}<16'b0011010101110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010101110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011010101110100) && ({row_reg, col_reg}<16'b0011010101110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010101110110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0011010101110111) && ({row_reg, col_reg}<16'b0011010101111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0011010101111011) && ({row_reg, col_reg}<16'b0011010101111101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0011010101111101) && ({row_reg, col_reg}<16'b0011010110000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011010110000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011010110000001) && ({row_reg, col_reg}<16'b0011010110000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010110000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011010110000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010110000101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011010110000110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011010110000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010110001000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0011010110001001) && ({row_reg, col_reg}<16'b0011010110001011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0011010110001011) && ({row_reg, col_reg}<16'b0011010110001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010110001110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011010110001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011010110010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010110010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011010110010010) && ({row_reg, col_reg}<16'b0011010110010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011010110010101) && ({row_reg, col_reg}<16'b0011010110010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011010110010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010110011000)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}==16'b0011010110011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010110011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011010110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011010110011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011010110011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011010110011111) && ({row_reg, col_reg}<16'b0011010110100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010110100011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011010110100100) && ({row_reg, col_reg}<16'b0011010110100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011010110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011010110101001) && ({row_reg, col_reg}<16'b0011010110101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011010110101100) && ({row_reg, col_reg}<16'b0011010110101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011010110101110) && ({row_reg, col_reg}<16'b0011010110110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011010110110000) && ({row_reg, col_reg}<16'b0011010110110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010110110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011010110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010110110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011010110110111) && ({row_reg, col_reg}<16'b0011010110111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010110111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011010110111010) && ({row_reg, col_reg}<16'b0011010110111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010110111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010110111101) && ({row_reg, col_reg}<16'b0011010111000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011010111000000) && ({row_reg, col_reg}<16'b0011010111000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011010111000101) && ({row_reg, col_reg}<16'b0011010111000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010111000111) && ({row_reg, col_reg}<16'b0011010111001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010111001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010111001011) && ({row_reg, col_reg}<16'b0011010111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010111010001) && ({row_reg, col_reg}<16'b0011010111101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011010111101111) && ({row_reg, col_reg}<16'b0011010111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010111110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010111110011) && ({row_reg, col_reg}<16'b0011010111110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010111110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011010111110111) && ({row_reg, col_reg}<16'b0011010111111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011010111111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010111111011) && ({row_reg, col_reg}<16'b0011010111111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0011010111111110) && ({row_reg, col_reg}<16'b0011011000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011000000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011011000000001) && ({row_reg, col_reg}<16'b0011011000000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011000000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011011000000100) && ({row_reg, col_reg}<16'b0011011000001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011000001000) && ({row_reg, col_reg}<16'b0011011000001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011011000001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011000001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011011000001100) && ({row_reg, col_reg}<16'b0011011000001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011000001110) && ({row_reg, col_reg}<16'b0011011000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011000010011) && ({row_reg, col_reg}<16'b0011011000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011011000100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011000100110) && ({row_reg, col_reg}<16'b0011011000101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011000101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011000101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011000101100) && ({row_reg, col_reg}<16'b0011011000101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011011000101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011011000101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011000110000) && ({row_reg, col_reg}<16'b0011011000110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011000110010) && ({row_reg, col_reg}<16'b0011011000110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011000110100) && ({row_reg, col_reg}<16'b0011011000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011011000110110) && ({row_reg, col_reg}<16'b0011011000111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011011000111001) && ({row_reg, col_reg}<16'b0011011000111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011000111100) && ({row_reg, col_reg}<16'b0011011000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011011000111110) && ({row_reg, col_reg}<16'b0011011001000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011001000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011011001000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011011001000101) && ({row_reg, col_reg}<16'b0011011001000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011011001000111) && ({row_reg, col_reg}<16'b0011011001001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011011001001100) && ({row_reg, col_reg}<16'b0011011001001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011011001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011011001001111) && ({row_reg, col_reg}<16'b0011011001010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011011001010010) && ({row_reg, col_reg}<16'b0011011001010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011001010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011011001010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011011001010111) && ({row_reg, col_reg}<16'b0011011001011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011001011001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011011001011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011011001011011) && ({row_reg, col_reg}<16'b0011011001011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011001100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011011001100001) && ({row_reg, col_reg}<16'b0011011001100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011011001100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011011001100101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011011001100110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011011001100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011011001101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011011001101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011011001101010)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0011011001101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011011001101100) && ({row_reg, col_reg}<16'b0011011001101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011011001101111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011011001110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011001110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011001110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011001110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011011001110100) && ({row_reg, col_reg}<16'b0011011001110111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0011011001110111) && ({row_reg, col_reg}<16'b0011011001111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0011011001111011) && ({row_reg, col_reg}<16'b0011011001111101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0011011001111101) && ({row_reg, col_reg}<16'b0011011010000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011011010000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011011010000001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011011010000010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011011010000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011011010000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011011010000101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011011010000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011011010000111) && ({row_reg, col_reg}<16'b0011011010001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011010001001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011011010001010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011011010001011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0011011010001100) && ({row_reg, col_reg}<16'b0011011010001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011011010001111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011011010010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011010010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011010010010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011011010010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011011010010100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0011011010010101) && ({row_reg, col_reg}<16'b0011011010010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011011010010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011010011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011010011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011011010011011) && ({row_reg, col_reg}<16'b0011011010011101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011011010011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011011010011110) && ({row_reg, col_reg}<16'b0011011010100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011011010100000) && ({row_reg, col_reg}<16'b0011011010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011010100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011011010100100) && ({row_reg, col_reg}<16'b0011011010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011011010100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011011010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011011010101001) && ({row_reg, col_reg}<16'b0011011010101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011011010101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011011010101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011011010101110) && ({row_reg, col_reg}<16'b0011011010110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011011010110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011011010110001)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011011010110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011011010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011010110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011011010110111) && ({row_reg, col_reg}<16'b0011011010111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011010111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011011010111010) && ({row_reg, col_reg}<16'b0011011010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011010111101) && ({row_reg, col_reg}<16'b0011011011000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011011011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011011000001) && ({row_reg, col_reg}<16'b0011011011000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011011011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011011011000100) && ({row_reg, col_reg}<16'b0011011011000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011011000111) && ({row_reg, col_reg}<16'b0011011011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011011001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011011001011) && ({row_reg, col_reg}<16'b0011011011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011011010001) && ({row_reg, col_reg}<16'b0011011011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011011011101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011011110000) && ({row_reg, col_reg}<16'b0011011011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011011110010) && ({row_reg, col_reg}<16'b0011011011110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011011011110110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=16'b0011011011110111) && ({row_reg, col_reg}<16'b0011011011111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011011111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011011011111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011011111011) && ({row_reg, col_reg}<16'b0011011011111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0011011011111110) && ({row_reg, col_reg}<16'b0011011100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011100000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011011100000001) && ({row_reg, col_reg}<16'b0011011100000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011100000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011011100000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011100000101) && ({row_reg, col_reg}<16'b0011011100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011011100001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011011100001001) && ({row_reg, col_reg}<16'b0011011100001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011100001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011011100001100) && ({row_reg, col_reg}<16'b0011011100001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011100001110) && ({row_reg, col_reg}<16'b0011011100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011100010011) && ({row_reg, col_reg}<16'b0011011100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011011100100110) && ({row_reg, col_reg}<16'b0011011100101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011100101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011100101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011100101100) && ({row_reg, col_reg}<16'b0011011100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011011100101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011011100101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011100110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011100110001) && ({row_reg, col_reg}<16'b0011011100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011011100110011) && ({row_reg, col_reg}<16'b0011011100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011100110110) && ({row_reg, col_reg}<16'b0011011100111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011100111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011100111010) && ({row_reg, col_reg}<16'b0011011100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011100111110) && ({row_reg, col_reg}<16'b0011011101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011101000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011011101000100) && ({row_reg, col_reg}<16'b0011011101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011011101000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011101001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011101001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011011101001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011011101001011) && ({row_reg, col_reg}<16'b0011011101001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011011101001101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011011101001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011011101001111) && ({row_reg, col_reg}<16'b0011011101010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011011101010010) && ({row_reg, col_reg}<16'b0011011101010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011101010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011101010110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011011101010111) && ({row_reg, col_reg}<16'b0011011101011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011011101011001) && ({row_reg, col_reg}<16'b0011011101011011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011011101011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011011101011100) && ({row_reg, col_reg}<16'b0011011101011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011101011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011101100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011011101100001) && ({row_reg, col_reg}<16'b0011011101100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011011101100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011011101100101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011011101100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011101100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011011101101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011011101101001) && ({row_reg, col_reg}<16'b0011011101101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011101101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011011101101100) && ({row_reg, col_reg}<16'b0011011101101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011011101101111) && ({row_reg, col_reg}<16'b0011011101110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011101110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011011101110011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011011101110100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0011011101110101) && ({row_reg, col_reg}<16'b0011011101110111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0011011101110111) && ({row_reg, col_reg}<16'b0011011101111001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011011101111001)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011011101111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011011101111011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011011101111100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0011011101111101) && ({row_reg, col_reg}<16'b0011011101111111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011011101111111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0011011110000000) && ({row_reg, col_reg}<16'b0011011110000010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011011110000010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011011110000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011011110000100) && ({row_reg, col_reg}<16'b0011011110000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011011110000111) && ({row_reg, col_reg}<16'b0011011110001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011110001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011011110001010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0011011110001011) && ({row_reg, col_reg}<16'b0011011110001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011011110001111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011011110010000) && ({row_reg, col_reg}<16'b0011011110010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011011110010010) && ({row_reg, col_reg}<16'b0011011110010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011011110010101) && ({row_reg, col_reg}<16'b0011011110010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011011110010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011110011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011110011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011011110011011) && ({row_reg, col_reg}<16'b0011011110011101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011011110011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011011110011110) && ({row_reg, col_reg}<16'b0011011110100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011011110100000) && ({row_reg, col_reg}<16'b0011011110100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011011110100011) && ({row_reg, col_reg}<16'b0011011110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011011110100110) && ({row_reg, col_reg}<16'b0011011110101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011011110101001) && ({row_reg, col_reg}<16'b0011011110101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011011110101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011011110101100) && ({row_reg, col_reg}<16'b0011011110101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011110101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011011110101111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011011110110000) && ({row_reg, col_reg}<16'b0011011110110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011011110110010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011011110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011110110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011011110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011110110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011011110110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011011110111001) && ({row_reg, col_reg}<16'b0011011110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011110111101) && ({row_reg, col_reg}<16'b0011011111000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011011111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011111000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011111000010) && ({row_reg, col_reg}<16'b0011011111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011011111000100) && ({row_reg, col_reg}<16'b0011011111000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011111000111) && ({row_reg, col_reg}<16'b0011011111001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011111001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011011111001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011111001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011011111001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011011111001111) && ({row_reg, col_reg}<16'b0011011111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011111010001) && ({row_reg, col_reg}<16'b0011011111110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011011111110000) && ({row_reg, col_reg}<16'b0011011111110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011111110010) && ({row_reg, col_reg}<16'b0011011111110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011111110111) && ({row_reg, col_reg}<16'b0011011111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011011111111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011011111111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011111111011) && ({row_reg, col_reg}<16'b0011011111111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0011011111111110) && ({row_reg, col_reg}<16'b0011100000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100000000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011100000000001) && ({row_reg, col_reg}<16'b0011100000000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011100000000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011100000000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100000000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011100000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100000000111) && ({row_reg, col_reg}<16'b0011100000001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011100000001001) && ({row_reg, col_reg}<16'b0011100000001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011100000001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011100000001100) && ({row_reg, col_reg}<16'b0011100000001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100000001110) && ({row_reg, col_reg}<16'b0011100000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100000010011) && ({row_reg, col_reg}<16'b0011100000100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011100000100110) && ({row_reg, col_reg}<16'b0011100000101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100000101000) && ({row_reg, col_reg}<16'b0011100000101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100000101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011100000101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011100000101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100000101110) && ({row_reg, col_reg}<16'b0011100000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100000110000) && ({row_reg, col_reg}<16'b0011100000110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011100000110011) && ({row_reg, col_reg}<16'b0011100000110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100000110110) && ({row_reg, col_reg}<16'b0011100000111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100000111001) && ({row_reg, col_reg}<16'b0011100000111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100000111111) && ({row_reg, col_reg}<16'b0011100001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100001000001) && ({row_reg, col_reg}<16'b0011100001000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011100001000100) && ({row_reg, col_reg}<16'b0011100001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011100001000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011100001000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100001001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100001001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011100001001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100001001011) && ({row_reg, col_reg}<16'b0011100001001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011100001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100001001111) && ({row_reg, col_reg}<16'b0011100001010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011100001010010) && ({row_reg, col_reg}<16'b0011100001010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100001010101) && ({row_reg, col_reg}<16'b0011100001011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100001011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011100001011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011100001011011) && ({row_reg, col_reg}<16'b0011100001011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011100001011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100001011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011100001100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011100001100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011100001100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011100001100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011100001100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011100001100101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011100001100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100001100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011100001101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011100001101001) && ({row_reg, col_reg}<16'b0011100001101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011100001101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011100001101100) && ({row_reg, col_reg}<16'b0011100001101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011100001101110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011100001101111) && ({row_reg, col_reg}<16'b0011100001110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100001110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011100001110010) && ({row_reg, col_reg}<16'b0011100001110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0011100001110101) && ({row_reg, col_reg}<16'b0011100001111000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011100001111000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011100001111001)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}>=16'b0011100001111010) && ({row_reg, col_reg}<16'b0011100001111100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011100001111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011100001111101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011100001111110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011100001111111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0011100010000000) && ({row_reg, col_reg}<16'b0011100010000010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011100010000010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011100010000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011100010000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011100010000101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011100010000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011100010000111) && ({row_reg, col_reg}<16'b0011100010001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100010001001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011100010001010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011100010001011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011100010001100) && ({row_reg, col_reg}<16'b0011100010001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011100010001110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011100010001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011100010010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100010010001) && ({row_reg, col_reg}<16'b0011100010010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100010010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011100010010100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0011100010010101) && ({row_reg, col_reg}<16'b0011100010010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011100010010111) && ({row_reg, col_reg}<16'b0011100010011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011100010011011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011100010011100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011100010011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011100010011110) && ({row_reg, col_reg}<16'b0011100010100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100010100000) && ({row_reg, col_reg}<16'b0011100010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011100010100011) && ({row_reg, col_reg}<16'b0011100010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011100010100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011100010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100010101001) && ({row_reg, col_reg}<16'b0011100010101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011100010101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011100010101100) && ({row_reg, col_reg}<16'b0011100010101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011100010101110) && ({row_reg, col_reg}<16'b0011100010110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100010110000) && ({row_reg, col_reg}<16'b0011100010110011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011100010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100010110101) && ({row_reg, col_reg}<16'b0011100010110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011100010110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011100010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011100010111001) && ({row_reg, col_reg}<16'b0011100010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100010111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100010111110) && ({row_reg, col_reg}<16'b0011100011000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011100011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100011000010) && ({row_reg, col_reg}<16'b0011100011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011100011000100) && ({row_reg, col_reg}<16'b0011100011001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011100011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100011001001) && ({row_reg, col_reg}<16'b0011100011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100011001011) && ({row_reg, col_reg}<16'b0011100011001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100011001111) && ({row_reg, col_reg}<16'b0011100011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100011010001) && ({row_reg, col_reg}<16'b0011100011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011100011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100011110000) && ({row_reg, col_reg}<16'b0011100011110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100011110010) && ({row_reg, col_reg}<16'b0011100011110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100011110100) && ({row_reg, col_reg}<16'b0011100011110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100011110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100011110111) && ({row_reg, col_reg}<16'b0011100011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011100011111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011100011111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100011111011) && ({row_reg, col_reg}<16'b0011100011111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0011100011111110) && ({row_reg, col_reg}<16'b0011100100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100100000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011100100000001) && ({row_reg, col_reg}<16'b0011100100000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011100100000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011100100000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100100000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011100100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100100000111) && ({row_reg, col_reg}<16'b0011100100001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011100100001001) && ({row_reg, col_reg}<16'b0011100100001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011100100001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011100100001100) && ({row_reg, col_reg}<16'b0011100100001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100100001110) && ({row_reg, col_reg}<16'b0011100100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100100010011) && ({row_reg, col_reg}<16'b0011100100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011100100100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100100100110) && ({row_reg, col_reg}<16'b0011100100101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100100101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011100100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011100100101101) && ({row_reg, col_reg}<16'b0011100100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100100110000) && ({row_reg, col_reg}<16'b0011100100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011100100110010) && ({row_reg, col_reg}<16'b0011100100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100100110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011100100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100100110110) && ({row_reg, col_reg}<16'b0011100100111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100100111001) && ({row_reg, col_reg}<16'b0011100100111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100100111100) && ({row_reg, col_reg}<16'b0011100100111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011100100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100100111111) && ({row_reg, col_reg}<16'b0011100101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100101000001) && ({row_reg, col_reg}<16'b0011100101000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011100101000100) && ({row_reg, col_reg}<16'b0011100101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011100101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011100101000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100101001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100101001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011100101001010) && ({row_reg, col_reg}<16'b0011100101001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011100101001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011100101001101) && ({row_reg, col_reg}<16'b0011100101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100101001111) && ({row_reg, col_reg}<16'b0011100101010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011100101010011) && ({row_reg, col_reg}<16'b0011100101010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011100101010101) && ({row_reg, col_reg}<16'b0011100101011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011100101011001) && ({row_reg, col_reg}<16'b0011100101011011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011100101011011) && ({row_reg, col_reg}<16'b0011100101011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011100101011111) && ({row_reg, col_reg}<16'b0011100101100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011100101100001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0011100101100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011100101100011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0011100101100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011100101100101) && ({row_reg, col_reg}<16'b0011100101100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100101100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011100101101000) && ({row_reg, col_reg}<16'b0011100101101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011100101101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011100101101100) && ({row_reg, col_reg}<16'b0011100101101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011100101101110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011100101101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100101110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011100101110001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011100101110010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0011100101110011) && ({row_reg, col_reg}<16'b0011100101110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011100101110111)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0011100101111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011100101111001)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011100101111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011100101111011)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0011100101111100) && ({row_reg, col_reg}<16'b0011100101111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011100101111110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011100101111111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011100110000000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011100110000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011100110000010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011100110000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011100110000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011100110000101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011100110000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011100110000111) && ({row_reg, col_reg}<16'b0011100110001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100110001001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011100110001010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011100110001011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011100110001100) && ({row_reg, col_reg}<16'b0011100110001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011100110001110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011100110001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011100110010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011100110010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011100110010010) && ({row_reg, col_reg}<16'b0011100110010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011100110010100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0011100110010101) && ({row_reg, col_reg}<16'b0011100110010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011100110010111) && ({row_reg, col_reg}<16'b0011100110011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011100110011011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011100110011100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011100110011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011100110011110) && ({row_reg, col_reg}<16'b0011100110100100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011100110100100) && ({row_reg, col_reg}<16'b0011100110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011100110100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011100110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100110101001) && ({row_reg, col_reg}<16'b0011100110101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011100110101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011100110101100) && ({row_reg, col_reg}<16'b0011100110101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011100110101110) && ({row_reg, col_reg}<16'b0011100110110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011100110110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011100110110001) && ({row_reg, col_reg}<16'b0011100110110100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011100110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100110110101) && ({row_reg, col_reg}<16'b0011100110111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011100110111001) && ({row_reg, col_reg}<16'b0011100110111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100110111111) && ({row_reg, col_reg}<16'b0011100111000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011100111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100111000010) && ({row_reg, col_reg}<16'b0011100111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011100111000100) && ({row_reg, col_reg}<16'b0011100111001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011100111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100111001001) && ({row_reg, col_reg}<16'b0011100111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100111001011) && ({row_reg, col_reg}<16'b0011100111001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100111001101) && ({row_reg, col_reg}<16'b0011100111001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011100111001111) && ({row_reg, col_reg}<16'b0011100111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100111010001) && ({row_reg, col_reg}<16'b0011100111101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011100111101111) && ({row_reg, col_reg}<16'b0011100111110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100111110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100111110011) && ({row_reg, col_reg}<16'b0011100111110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100111110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100111110111) && ({row_reg, col_reg}<16'b0011100111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011100111111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011100111111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100111111011) && ({row_reg, col_reg}<16'b0011100111111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011100111111110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}==16'b0011100111111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011101000000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011101000000001) && ({row_reg, col_reg}<16'b0011101000000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101000000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011101000000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101000000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011101000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101000000111) && ({row_reg, col_reg}<16'b0011101000001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011101000001001) && ({row_reg, col_reg}<16'b0011101000001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101000001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011101000001100) && ({row_reg, col_reg}<16'b0011101000001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101000001110) && ({row_reg, col_reg}<16'b0011101000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011101000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101000010011) && ({row_reg, col_reg}<16'b0011101000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011101000100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101000100110) && ({row_reg, col_reg}<16'b0011101000101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101000101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011101000101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011101000101101) && ({row_reg, col_reg}<16'b0011101000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101000110000) && ({row_reg, col_reg}<16'b0011101000110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101000110010) && ({row_reg, col_reg}<16'b0011101000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101000110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011101000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101000110110) && ({row_reg, col_reg}<16'b0011101000111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101000111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011101000111010) && ({row_reg, col_reg}<16'b0011101000111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101000111100) && ({row_reg, col_reg}<16'b0011101000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011101000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101000111111) && ({row_reg, col_reg}<16'b0011101001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011101001000001) && ({row_reg, col_reg}<16'b0011101001000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011101001000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101001000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011101001000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101001001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011101001001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011101001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011101001001011) && ({row_reg, col_reg}<16'b0011101001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101001001111) && ({row_reg, col_reg}<16'b0011101001010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101001010010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011101001010011) && ({row_reg, col_reg}<16'b0011101001010101)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}>=16'b0011101001010101) && ({row_reg, col_reg}<16'b0011101001011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011101001011001) && ({row_reg, col_reg}<16'b0011101001011011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011101001011011) && ({row_reg, col_reg}<16'b0011101001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101001011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011101001100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011101001100001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0011101001100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011101001100011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0011101001100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011101001100101) && ({row_reg, col_reg}<16'b0011101001100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101001100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011101001101000) && ({row_reg, col_reg}<16'b0011101001101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101001101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101001101011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011101001101100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011101001101101) && ({row_reg, col_reg}<16'b0011101001101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011101001101111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011101001110000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011101001110001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011101001110010)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0011101001110011) && ({row_reg, col_reg}<16'b0011101001110101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011101001110101) && ({row_reg, col_reg}<16'b0011101001110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011101001110111) && ({row_reg, col_reg}<16'b0011101001111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011101001111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0011101001111100) && ({row_reg, col_reg}<16'b0011101001111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011101001111110) && ({row_reg, col_reg}<16'b0011101010000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011101010000000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011101010000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011101010000010) && ({row_reg, col_reg}<16'b0011101010000100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011101010000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011101010000101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011101010000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011101010000111) && ({row_reg, col_reg}<16'b0011101010001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101010001001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011101010001010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011101010001011) && ({row_reg, col_reg}<16'b0011101010001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011101010001101) && ({row_reg, col_reg}<16'b0011101010001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011101010001111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011101010010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101010010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011101010010010) && ({row_reg, col_reg}<16'b0011101010010101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011101010010101) && ({row_reg, col_reg}<16'b0011101010010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011101010010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101010011000) && ({row_reg, col_reg}<16'b0011101010011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011101010011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011101010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011101010011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011101010011110) && ({row_reg, col_reg}<16'b0011101010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101010100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101010100100) && ({row_reg, col_reg}<16'b0011101010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011101010100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011101010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101010101001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0011101010101010) && ({row_reg, col_reg}<16'b0011101010110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101010110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011101010110001) && ({row_reg, col_reg}<16'b0011101010110011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011101010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101010110101) && ({row_reg, col_reg}<16'b0011101010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011101010111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011101010111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101010111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011101010111011) && ({row_reg, col_reg}<16'b0011101010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011101010111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011101011000000) && ({row_reg, col_reg}<16'b0011101011000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101011000010) && ({row_reg, col_reg}<16'b0011101011001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011101011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101011001001) && ({row_reg, col_reg}<16'b0011101011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011101011001011) && ({row_reg, col_reg}<16'b0011101011001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101011001101) && ({row_reg, col_reg}<16'b0011101011001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011101011001111) && ({row_reg, col_reg}<16'b0011101011010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101011010001) && ({row_reg, col_reg}<16'b0011101011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011101011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101011110000) && ({row_reg, col_reg}<16'b0011101011110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011101011110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101011110011) && ({row_reg, col_reg}<16'b0011101011110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101011110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011101011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011101011111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011101011111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101011111011) && ({row_reg, col_reg}<16'b0011101011111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0011101011111110) && ({row_reg, col_reg}<16'b0011101100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101100000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011101100000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101100000010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0011101100000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011101100000100) && ({row_reg, col_reg}<16'b0011101100001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011101100001001) && ({row_reg, col_reg}<16'b0011101100001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101100001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011101100001100) && ({row_reg, col_reg}<16'b0011101100001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101100001110) && ({row_reg, col_reg}<16'b0011101100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011101100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101100010011) && ({row_reg, col_reg}<16'b0011101100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011101100100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101100100110) && ({row_reg, col_reg}<16'b0011101100101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101100101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011101100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011101100101101) && ({row_reg, col_reg}<16'b0011101100110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101100110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101100110010) && ({row_reg, col_reg}<16'b0011101100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101100110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011101100110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011101100110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011101100110111) && ({row_reg, col_reg}<16'b0011101100111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101100111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011101100111010) && ({row_reg, col_reg}<16'b0011101100111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101100111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011101100111101) && ({row_reg, col_reg}<16'b0011101100111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101100111111) && ({row_reg, col_reg}<16'b0011101101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011101101000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011101101000010) && ({row_reg, col_reg}<16'b0011101101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011101101000111) && ({row_reg, col_reg}<16'b0011101101001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011101101001001) && ({row_reg, col_reg}<16'b0011101101001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101101001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011101101001101) && ({row_reg, col_reg}<16'b0011101101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101101001111) && ({row_reg, col_reg}<16'b0011101101010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011101101010010) && ({row_reg, col_reg}<16'b0011101101010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011101101010101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011101101010110) && ({row_reg, col_reg}<16'b0011101101011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011101101011001) && ({row_reg, col_reg}<16'b0011101101011011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011101101011011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011101101011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011101101011101) && ({row_reg, col_reg}<16'b0011101101100000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011101101100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011101101100001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0011101101100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011101101100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011101101100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011101101100101) && ({row_reg, col_reg}<16'b0011101101100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101101100111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011101101101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011101101101001) && ({row_reg, col_reg}<16'b0011101101101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101101101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011101101101100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011101101101101) && ({row_reg, col_reg}<16'b0011101101101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011101101101111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011101101110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011101101110001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011101101110010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011101101110011)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0011101101110100) && ({row_reg, col_reg}<16'b0011101101110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011101101110111) && ({row_reg, col_reg}<16'b0011101101111001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011101101111001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0011101101111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0011101101111011) && ({row_reg, col_reg}<16'b0011101101111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011101101111101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011101101111110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011101101111111)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0011101110000000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011101110000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011101110000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101110000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011101110000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011101110000101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011101110000110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011101110000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011101110001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101110001001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0011101110001010) && ({row_reg, col_reg}<16'b0011101110001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011101110001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011101110001110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011101110001111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0011101110010000) && ({row_reg, col_reg}<16'b0011101110010010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011101110010010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0011101110010011) && ({row_reg, col_reg}<16'b0011101110010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101110010101)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011101110010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011101110010111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011101110011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101110011001)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011101110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011101110011011) && ({row_reg, col_reg}<16'b0011101110011101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011101110011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011101110011110) && ({row_reg, col_reg}<16'b0011101110100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101110100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011101110100001) && ({row_reg, col_reg}<16'b0011101110100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101110100100) && ({row_reg, col_reg}<16'b0011101110100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011101110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011101110101000) && ({row_reg, col_reg}<16'b0011101110101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101110101101) && ({row_reg, col_reg}<16'b0011101110110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101110110001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011101110110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011101110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101110110101) && ({row_reg, col_reg}<16'b0011101110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011101110111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011101110111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101110111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011101110111011) && ({row_reg, col_reg}<16'b0011101110111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011101110111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011101111000000) && ({row_reg, col_reg}<16'b0011101111000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101111000010) && ({row_reg, col_reg}<16'b0011101111000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101111000111) && ({row_reg, col_reg}<16'b0011101111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101111001001) && ({row_reg, col_reg}<16'b0011101111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011101111001011) && ({row_reg, col_reg}<16'b0011101111001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101111001101) && ({row_reg, col_reg}<16'b0011101111001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011101111001111) && ({row_reg, col_reg}<16'b0011101111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101111010001) && ({row_reg, col_reg}<16'b0011101111110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011101111110000) && ({row_reg, col_reg}<16'b0011101111110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011101111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101111110011) && ({row_reg, col_reg}<16'b0011101111110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011101111110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101111110111) && ({row_reg, col_reg}<16'b0011101111111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011101111111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101111111011) && ({row_reg, col_reg}<16'b0011101111111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0011101111111110) && ({row_reg, col_reg}<16'b0011110000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110000000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011110000000001) && ({row_reg, col_reg}<16'b0011110000000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011110000000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011110000000100) && ({row_reg, col_reg}<16'b0011110000001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110000001000) && ({row_reg, col_reg}<16'b0011110000001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011110000001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011110000001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110000001100) && ({row_reg, col_reg}<16'b0011110000001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110000001110) && ({row_reg, col_reg}<16'b0011110000010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110000010011) && ({row_reg, col_reg}<16'b0011110000100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011110000100110) && ({row_reg, col_reg}<16'b0011110000101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110000101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011110000101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011110000101101) && ({row_reg, col_reg}<16'b0011110000110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110000110011) && ({row_reg, col_reg}<16'b0011110000110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011110000110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011110000111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011110000111001) && ({row_reg, col_reg}<16'b0011110001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110001000001) && ({row_reg, col_reg}<16'b0011110001000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011110001000011) && ({row_reg, col_reg}<16'b0011110001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011110001000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011110001000111) && ({row_reg, col_reg}<16'b0011110001001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110001001001) && ({row_reg, col_reg}<16'b0011110001001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110001001100) && ({row_reg, col_reg}<16'b0011110001001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011110001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110001001111) && ({row_reg, col_reg}<16'b0011110001010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110001010010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011110001010011)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0011110001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011110001010101) && ({row_reg, col_reg}<16'b0011110001011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011110001011000) && ({row_reg, col_reg}<16'b0011110001011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011110001011100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011110001011101) && ({row_reg, col_reg}<16'b0011110001100000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011110001100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011110001100001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0011110001100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011110001100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011110001100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011110001100101) && ({row_reg, col_reg}<16'b0011110001100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110001100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011110001101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011110001101001) && ({row_reg, col_reg}<16'b0011110001101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011110001101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011110001101100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011110001101101) && ({row_reg, col_reg}<16'b0011110001101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011110001101111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011110001110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011110001110001) && ({row_reg, col_reg}<16'b0011110001110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011110001110011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011110001110100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011110001110101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011110001110110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011110001110111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011110001111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011110001111001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0011110001111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011110001111011)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0011110001111100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0011110001111101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011110001111110)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011110001111111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011110010000000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011110010000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011110010000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110010000011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011110010000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011110010000101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011110010000110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011110010000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011110010001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110010001001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0011110010001010) && ({row_reg, col_reg}<16'b0011110010001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011110010001101) && ({row_reg, col_reg}<16'b0011110010010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110010010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011110010010001) && ({row_reg, col_reg}<16'b0011110010010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011110010010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110010010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110010010101) && ({row_reg, col_reg}<16'b0011110010011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011110010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011110010011011) && ({row_reg, col_reg}<16'b0011110010011101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011110010011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011110010011110) && ({row_reg, col_reg}<16'b0011110010100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011110010100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011110010100011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011110010100100) && ({row_reg, col_reg}<16'b0011110010100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011110010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011110010101000) && ({row_reg, col_reg}<16'b0011110010101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110010101011) && ({row_reg, col_reg}<16'b0011110010110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110010110001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011110010110010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011110010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110010110101) && ({row_reg, col_reg}<16'b0011110010110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110010110111) && ({row_reg, col_reg}<16'b0011110010111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011110010111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011110010111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011110010111011) && ({row_reg, col_reg}<16'b0011110010111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110010111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011110010111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011110011000000) && ({row_reg, col_reg}<16'b0011110011000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110011000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011110011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011110011000100) && ({row_reg, col_reg}<16'b0011110011000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110011000111) && ({row_reg, col_reg}<16'b0011110011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110011001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011110011001100) && ({row_reg, col_reg}<16'b0011110011001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110011001111) && ({row_reg, col_reg}<16'b0011110011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110011010001) && ({row_reg, col_reg}<16'b0011110011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011110011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110011110001) && ({row_reg, col_reg}<16'b0011110011110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110011110011) && ({row_reg, col_reg}<16'b0011110011110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110011110110) && ({row_reg, col_reg}<16'b0011110011111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110011111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110011111011) && ({row_reg, col_reg}<16'b0011110011111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0011110011111110) && ({row_reg, col_reg}<16'b0011110100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110100000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011110100000001) && ({row_reg, col_reg}<16'b0011110100000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011110100000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011110100000101) && ({row_reg, col_reg}<16'b0011110100000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110100001000) && ({row_reg, col_reg}<16'b0011110100001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011110100001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011110100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110100001100) && ({row_reg, col_reg}<16'b0011110100001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110100001110) && ({row_reg, col_reg}<16'b0011110100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110100010011) && ({row_reg, col_reg}<16'b0011110100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011110100100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110100100111) && ({row_reg, col_reg}<16'b0011110100101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110100101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011110100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011110100101101) && ({row_reg, col_reg}<16'b0011110100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110100110100) && ({row_reg, col_reg}<16'b0011110100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110100110110) && ({row_reg, col_reg}<16'b0011110100111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011110100111001) && ({row_reg, col_reg}<16'b0011110100111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110100111100) && ({row_reg, col_reg}<16'b0011110100111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011110100111110) && ({row_reg, col_reg}<16'b0011110101000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110101000010) && ({row_reg, col_reg}<16'b0011110101000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011110101000100) && ({row_reg, col_reg}<16'b0011110101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011110101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011110101000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110101001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110101001001) && ({row_reg, col_reg}<16'b0011110101001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110101001100) && ({row_reg, col_reg}<16'b0011110101001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011110101001110) && ({row_reg, col_reg}<16'b0011110101010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110101010010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011110101010011)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0011110101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011110101010101) && ({row_reg, col_reg}<16'b0011110101011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011110101011001) && ({row_reg, col_reg}<16'b0011110101011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011110101011100) && ({row_reg, col_reg}<16'b0011110101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110101011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011110101011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011110101100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011110101100001) && ({row_reg, col_reg}<16'b0011110101100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0011110101100100) && ({row_reg, col_reg}<16'b0011110101101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011110101101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110101101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011110101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110101101011) && ({row_reg, col_reg}<16'b0011110101101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011110101101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011110101101110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011110101101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110101110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011110101110001) && ({row_reg, col_reg}<16'b0011110101110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011110101110011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011110101110100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011110101110101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011110101110110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011110101110111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011110101111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011110101111001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0011110101111010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011110101111011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011110101111100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011110101111101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0011110101111110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011110101111111)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0011110110000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011110110000001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011110110000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110110000011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011110110000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011110110000101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011110110000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011110110000111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011110110001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110110001001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0011110110001010) && ({row_reg, col_reg}<16'b0011110110001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011110110001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011110110001110) && ({row_reg, col_reg}<16'b0011110110010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011110110010001) && ({row_reg, col_reg}<16'b0011110110010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011110110010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110110011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011110110011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011110110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011110110011011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011110110011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011110110011101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011110110011110) && ({row_reg, col_reg}<16'b0011110110100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011110110100000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011110110100001) && ({row_reg, col_reg}<16'b0011110110100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110110100011) && ({row_reg, col_reg}<16'b0011110110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011110110100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011110110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011110110101001) && ({row_reg, col_reg}<16'b0011110110101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110110101011) && ({row_reg, col_reg}<16'b0011110110110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011110110110000) && ({row_reg, col_reg}<16'b0011110110110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011110110110010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011110110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011110110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110110110110) && ({row_reg, col_reg}<16'b0011110110111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110110111001) && ({row_reg, col_reg}<16'b0011110110111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011110110111100) && ({row_reg, col_reg}<16'b0011110110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110110111110) && ({row_reg, col_reg}<16'b0011110111000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011110111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110111000010) && ({row_reg, col_reg}<16'b0011110111000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011110111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110111001000) && ({row_reg, col_reg}<16'b0011110111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110111001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011110111001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110111001101) && ({row_reg, col_reg}<16'b0011110111001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110111001111) && ({row_reg, col_reg}<16'b0011110111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110111010001) && ({row_reg, col_reg}<16'b0011110111101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011110111101111) && ({row_reg, col_reg}<16'b0011110111110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110111110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110111110101) && ({row_reg, col_reg}<16'b0011110111110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110111110111) && ({row_reg, col_reg}<16'b0011110111111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110111111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110111111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110111111011) && ({row_reg, col_reg}<16'b0011110111111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0011110111111110) && ({row_reg, col_reg}<16'b0011111000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111000000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011111000000001) && ({row_reg, col_reg}<16'b0011111000000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011111000000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111000000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011111000000101) && ({row_reg, col_reg}<16'b0011111000000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111000000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011111000001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011111000001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011111000001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111000001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011111000001100) && ({row_reg, col_reg}<16'b0011111000001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111000001110) && ({row_reg, col_reg}<16'b0011111000010000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011111000010000) && ({row_reg, col_reg}<16'b0011111000010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011111000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111000010011) && ({row_reg, col_reg}<16'b0011111000100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111000100111) && ({row_reg, col_reg}<16'b0011111000101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011111000101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011111000101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111000101101) && ({row_reg, col_reg}<16'b0011111000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111000110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111000110010) && ({row_reg, col_reg}<16'b0011111000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111000110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011111000110101) && ({row_reg, col_reg}<16'b0011111000110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111000110111) && ({row_reg, col_reg}<16'b0011111000111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011111000111001) && ({row_reg, col_reg}<16'b0011111000111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111000111100) && ({row_reg, col_reg}<16'b0011111000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011111000111110) && ({row_reg, col_reg}<16'b0011111001000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111001000100) && ({row_reg, col_reg}<16'b0011111001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111001000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011111001000111) && ({row_reg, col_reg}<16'b0011111001001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011111001001100) && ({row_reg, col_reg}<16'b0011111001001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011111001001110) && ({row_reg, col_reg}<16'b0011111001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111001010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011111001010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111001010010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011111001010011)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0011111001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011111001010101) && ({row_reg, col_reg}<16'b0011111001011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011111001011010) && ({row_reg, col_reg}<16'b0011111001011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011111001011101) && ({row_reg, col_reg}<16'b0011111001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111001011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111001100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011111001100001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011111001100010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011111001100011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0011111001100100) && ({row_reg, col_reg}<16'b0011111001101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011111001101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111001101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011111001101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011111001101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011111001101100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011111001101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011111001101110) && ({row_reg, col_reg}<16'b0011111001110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111001110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011111001110001) && ({row_reg, col_reg}<16'b0011111001110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011111001110011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011111001110100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011111001110101) && ({row_reg, col_reg}<16'b0011111001110111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011111001110111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011111001111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011111001111001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0011111001111010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011111001111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0011111001111100) && ({row_reg, col_reg}<16'b0011111001111111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111001111111)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0011111010000000) && ({row_reg, col_reg}<16'b0011111010000010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111010000010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011111010000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011111010000100) && ({row_reg, col_reg}<16'b0011111010000110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011111010000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011111010000111) && ({row_reg, col_reg}<16'b0011111010001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111010001001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0011111010001010) && ({row_reg, col_reg}<16'b0011111010001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011111010001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111010001110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011111010001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111010010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111010010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011111010010010) && ({row_reg, col_reg}<16'b0011111010010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011111010010111) && ({row_reg, col_reg}<16'b0011111010011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111010011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011111010011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011111010011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011111010011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011111010011110) && ({row_reg, col_reg}<16'b0011111010100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111010100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111010100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111010100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011111010100011) && ({row_reg, col_reg}<16'b0011111010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111010100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011111010100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011111010101001) && ({row_reg, col_reg}<16'b0011111010101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011111010101011) && ({row_reg, col_reg}<16'b0011111010101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011111010101101) && ({row_reg, col_reg}<16'b0011111010101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011111010101111) && ({row_reg, col_reg}<16'b0011111010110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011111010110001) && ({row_reg, col_reg}<16'b0011111010110011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011111010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111010110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011111010110101)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b0011111010110110) && ({row_reg, col_reg}<16'b0011111010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011111010111001) && ({row_reg, col_reg}<16'b0011111010111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011111010111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011111010111100) && ({row_reg, col_reg}<16'b0011111010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011111010111110) && ({row_reg, col_reg}<16'b0011111011000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011111011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111011000010) && ({row_reg, col_reg}<16'b0011111011000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111011000111) && ({row_reg, col_reg}<16'b0011111011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111011001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011111011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111011001011) && ({row_reg, col_reg}<16'b0011111011001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011111011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111011001111) && ({row_reg, col_reg}<16'b0011111011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111011010001) && ({row_reg, col_reg}<16'b0011111011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111011101111) && ({row_reg, col_reg}<16'b0011111011110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111011110111) && ({row_reg, col_reg}<16'b0011111011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011111011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011111011111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111011111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011111011111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011111011111101)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0011111011111110) && ({row_reg, col_reg}<16'b0011111100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111100000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011111100000001) && ({row_reg, col_reg}<16'b0011111100000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011111100000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011111100000100) && ({row_reg, col_reg}<16'b0011111100001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011111100001001) && ({row_reg, col_reg}<16'b0011111100001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111100001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011111100001100) && ({row_reg, col_reg}<16'b0011111100001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111100001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011111100001111) && ({row_reg, col_reg}<16'b0011111100010001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011111100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011111100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111100010011) && ({row_reg, col_reg}<16'b0011111100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111100100100) && ({row_reg, col_reg}<16'b0011111100100110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011111100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111100100111) && ({row_reg, col_reg}<16'b0011111100101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011111100101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011111100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111100101101) && ({row_reg, col_reg}<16'b0011111100110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111100110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111100110010) && ({row_reg, col_reg}<16'b0011111100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111100110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011111100110101) && ({row_reg, col_reg}<16'b0011111100110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011111100110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111100111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011111100111001) && ({row_reg, col_reg}<16'b0011111100111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111100111100) && ({row_reg, col_reg}<16'b0011111100111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011111100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111100111111) && ({row_reg, col_reg}<16'b0011111101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111101000100) && ({row_reg, col_reg}<16'b0011111101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011111101000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111101001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011111101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011111101001100) && ({row_reg, col_reg}<16'b0011111101001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011111101001110) && ({row_reg, col_reg}<16'b0011111101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111101010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011111101010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111101010010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011111101010011)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0011111101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011111101010101) && ({row_reg, col_reg}<16'b0011111101011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111101011011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011111101011100) && ({row_reg, col_reg}<16'b0011111101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111101011110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011111101011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111101100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011111101100001) && ({row_reg, col_reg}<16'b0011111101100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011111101100011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011111101100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011111101100101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011111101100110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011111101100111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011111101101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011111101101001) && ({row_reg, col_reg}<16'b0011111101101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111101101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011111101101100) && ({row_reg, col_reg}<16'b0011111101101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011111101101110) && ({row_reg, col_reg}<16'b0011111101110001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111101110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011111101110010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0011111101110011) && ({row_reg, col_reg}<16'b0011111101110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011111101110111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0011111101111000) && ({row_reg, col_reg}<16'b0011111101111100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011111101111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011111101111101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111101111110)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}>=16'b0011111101111111) && ({row_reg, col_reg}<16'b0011111110000001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011111110000001) && ({row_reg, col_reg}<16'b0011111110000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111110000011)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0011111110000100) && ({row_reg, col_reg}<16'b0011111110000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011111110000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011111110000111) && ({row_reg, col_reg}<16'b0011111110001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111110001001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011111110001010) && ({row_reg, col_reg}<16'b0011111110001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011111110001110) && ({row_reg, col_reg}<16'b0011111110010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011111110010000) && ({row_reg, col_reg}<16'b0011111110010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011111110010010) && ({row_reg, col_reg}<16'b0011111110010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111110010100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0011111110010101) && ({row_reg, col_reg}<16'b0011111110010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011111110010111) && ({row_reg, col_reg}<16'b0011111110011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111110011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011111110011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011111110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011111110011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011111110011110) && ({row_reg, col_reg}<16'b0011111110100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111110100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111110100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111110100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011111110100011) && ({row_reg, col_reg}<16'b0011111110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111110100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011111110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111110101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011111110101010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011111110101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011111110101100) && ({row_reg, col_reg}<16'b0011111110101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011111110101110) && ({row_reg, col_reg}<16'b0011111110110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011111110110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011111110110001) && ({row_reg, col_reg}<16'b0011111110110011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011111110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111110110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011111110110101)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b0011111110110110) && ({row_reg, col_reg}<16'b0011111110111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111110111100) && ({row_reg, col_reg}<16'b0011111110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011111110111111) && ({row_reg, col_reg}<16'b0011111111000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011111111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111111000010) && ({row_reg, col_reg}<16'b0011111111000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111111000111) && ({row_reg, col_reg}<16'b0011111111001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111111001010) && ({row_reg, col_reg}<16'b0011111111001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011111111001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111111001111) && ({row_reg, col_reg}<16'b0011111111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111111010001) && ({row_reg, col_reg}<16'b0011111111110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111111110000) && ({row_reg, col_reg}<16'b0011111111110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111111110010) && ({row_reg, col_reg}<16'b0011111111110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111111110100) && ({row_reg, col_reg}<16'b0011111111110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111111110111) && ({row_reg, col_reg}<16'b0011111111111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011111111111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111111111010) && ({row_reg, col_reg}<16'b0011111111111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111111111100) && ({row_reg, col_reg}<16'b0011111111111110)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0011111111111110) && ({row_reg, col_reg}<16'b0100000000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000000000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000000000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100000000000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000000000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100000000000100) && ({row_reg, col_reg}<16'b0100000000001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000000001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100000000001001) && ({row_reg, col_reg}<16'b0100000000001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000000001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100000000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000000001101) && ({row_reg, col_reg}<16'b0100000000001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100000000001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000000010000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100000000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100000000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000000010011) && ({row_reg, col_reg}<16'b0100000000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100000000100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100000000100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000000100111) && ({row_reg, col_reg}<16'b0100000000101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100000000101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000000101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000000101101) && ({row_reg, col_reg}<16'b0100000000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000000110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100000000110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000000110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100000000110100) && ({row_reg, col_reg}<16'b0100000000110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100000000110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100000000111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100000000111001) && ({row_reg, col_reg}<16'b0100000000111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000000111100) && ({row_reg, col_reg}<16'b0100000000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100000000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000000111111) && ({row_reg, col_reg}<16'b0100000001000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100000001000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100000001000101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0100000001000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100000001000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000001001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100000001001001) && ({row_reg, col_reg}<16'b0100000001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100000001001011) && ({row_reg, col_reg}<16'b0100000001001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100000001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100000001001111) && ({row_reg, col_reg}<16'b0100000001010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000001010001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100000001010010) && ({row_reg, col_reg}<16'b0100000001010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100000001010101) && ({row_reg, col_reg}<16'b0100000001010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100000001010111) && ({row_reg, col_reg}<16'b0100000001011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100000001011010) && ({row_reg, col_reg}<16'b0100000001011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100000001011100) && ({row_reg, col_reg}<16'b0100000001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000001011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100000001100000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0100000001100001) && ({row_reg, col_reg}<16'b0100000001100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100000001100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100000001100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000001100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000001100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100000001101000) && ({row_reg, col_reg}<16'b0100000001101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000001101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000001101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100000001101100) && ({row_reg, col_reg}<16'b0100000001101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100000001101111) && ({row_reg, col_reg}<16'b0100000001110001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000001110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100000001110010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0100000001110011) && ({row_reg, col_reg}<16'b0100000001110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100000001110110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100000001110111) && ({row_reg, col_reg}<16'b0100000001111001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0100000001111001) && ({row_reg, col_reg}<16'b0100000001111011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0100000001111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0100000001111100) && ({row_reg, col_reg}<16'b0100000001111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100000001111110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100000001111111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100000010000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100000010000001) && ({row_reg, col_reg}<16'b0100000010000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000010000011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100000010000100) && ({row_reg, col_reg}<16'b0100000010000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100000010000110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0100000010000111) && ({row_reg, col_reg}<16'b0100000010001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100000010001001) && ({row_reg, col_reg}<16'b0100000010001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100000010001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100000010010000) && ({row_reg, col_reg}<16'b0100000010010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100000010010010) && ({row_reg, col_reg}<16'b0100000010010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100000010010101) && ({row_reg, col_reg}<16'b0100000010010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100000010010111) && ({row_reg, col_reg}<16'b0100000010011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100000010011001) && ({row_reg, col_reg}<16'b0100000010011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100000010011011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100000010011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100000010011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100000010011110) && ({row_reg, col_reg}<16'b0100000010100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000010100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100000010100011) && ({row_reg, col_reg}<16'b0100000010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000010100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0100000010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000010101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100000010101010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000010101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100000010101100) && ({row_reg, col_reg}<16'b0100000010101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000010101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100000010101111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100000010110000) && ({row_reg, col_reg}<16'b0100000010110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000010110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100000010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100000010110101) && ({row_reg, col_reg}<16'b0100000010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100000010111101) && ({row_reg, col_reg}<16'b0100000011000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100000011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000011000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100000011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000011000100) && ({row_reg, col_reg}<16'b0100000011001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000011001000) && ({row_reg, col_reg}<16'b0100000011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000011001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000011001011) && ({row_reg, col_reg}<16'b0100000011001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100000011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000011001111) && ({row_reg, col_reg}<16'b0100000011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000011010001) && ({row_reg, col_reg}<16'b0100000011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000011110000) && ({row_reg, col_reg}<16'b0100000011110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100000011110011) && ({row_reg, col_reg}<16'b0100000011110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000011110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100000011111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000011111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100000011111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100000011111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000011111100) && ({row_reg, col_reg}<16'b0100000011111110)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0100000011111110) && ({row_reg, col_reg}<16'b0100000100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000100000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100000100000001) && ({row_reg, col_reg}<16'b0100000100000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000100000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100000100000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000100000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100000100000110) && ({row_reg, col_reg}<16'b0100000100001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100000100001001) && ({row_reg, col_reg}<16'b0100000100001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000100001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100000100001100) && ({row_reg, col_reg}<16'b0100000100001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000100001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100000100001111) && ({row_reg, col_reg}<16'b0100000100010001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100000100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100000100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000100010011) && ({row_reg, col_reg}<16'b0100000100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100000100100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000100100110) && ({row_reg, col_reg}<16'b0100000100101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000100101000) && ({row_reg, col_reg}<16'b0100000100101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100000100101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100000100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000100101101) && ({row_reg, col_reg}<16'b0100000100110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000100110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100000100110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100000100110100) && ({row_reg, col_reg}<16'b0100000100110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100000100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000100110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100000100111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100000100111001) && ({row_reg, col_reg}<16'b0100000100111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000100111100) && ({row_reg, col_reg}<16'b0100000100111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100000100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000100111111) && ({row_reg, col_reg}<16'b0100000101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100000101000001) && ({row_reg, col_reg}<16'b0100000101000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100000101000100) && ({row_reg, col_reg}<16'b0100000101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100000101000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000101001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100000101001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100000101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100000101001100) && ({row_reg, col_reg}<16'b0100000101001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100000101001110) && ({row_reg, col_reg}<16'b0100000101010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000101010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100000101010001) && ({row_reg, col_reg}<16'b0100000101010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000101010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100000101010110) && ({row_reg, col_reg}<16'b0100000101011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100000101011010) && ({row_reg, col_reg}<16'b0100000101011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100000101011100) && ({row_reg, col_reg}<16'b0100000101011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000101011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100000101100000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100000101100001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0100000101100010) && ({row_reg, col_reg}<16'b0100000101100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100000101100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100000101100101) && ({row_reg, col_reg}<16'b0100000101100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000101100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100000101101000) && ({row_reg, col_reg}<16'b0100000101101010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000101101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100000101101011) && ({row_reg, col_reg}<16'b0100000101101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100000101101101) && ({row_reg, col_reg}<16'b0100000101110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100000101110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000101110001)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0100000101110010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0100000101110011) && ({row_reg, col_reg}<16'b0100000101110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100000101110101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0100000101110110) && ({row_reg, col_reg}<16'b0100000101111000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100000101111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100000101111001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0100000101111010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100000101111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100000101111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100000101111101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100000101111110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0100000101111111) && ({row_reg, col_reg}<16'b0100000110000001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100000110000001) && ({row_reg, col_reg}<16'b0100000110000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000110000011)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0100000110000100) && ({row_reg, col_reg}<16'b0100000110000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100000110000110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100000110000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100000110001000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100000110001001) && ({row_reg, col_reg}<16'b0100000110001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100000110001011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100000110001100) && ({row_reg, col_reg}<16'b0100000110001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100000110001111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100000110010000) && ({row_reg, col_reg}<16'b0100000110010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000110010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000110010011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0100000110010100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0100000110010101) && ({row_reg, col_reg}<16'b0100000110010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000110010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000110011000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100000110011001) && ({row_reg, col_reg}<16'b0100000110011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100000110011101) && ({row_reg, col_reg}<16'b0100000110011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000110011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100000110100000) && ({row_reg, col_reg}<16'b0100000110100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100000110100011) && ({row_reg, col_reg}<16'b0100000110100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100000110100111) && ({row_reg, col_reg}<16'b0100000110101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000110101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000110101010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000110101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100000110101100) && ({row_reg, col_reg}<16'b0100000110101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000110101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000110110000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0100000110110001) && ({row_reg, col_reg}<16'b0100000110110011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000110110011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100000110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100000110110101) && ({row_reg, col_reg}<16'b0100000110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100000110111101) && ({row_reg, col_reg}<16'b0100000111000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100000111000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100000111000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100000111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000111000100) && ({row_reg, col_reg}<16'b0100000111000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000111000111) && ({row_reg, col_reg}<16'b0100000111001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000111001010) && ({row_reg, col_reg}<16'b0100000111001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000111001111) && ({row_reg, col_reg}<16'b0100000111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000111010001) && ({row_reg, col_reg}<16'b0100000111110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100000111110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000111110001) && ({row_reg, col_reg}<16'b0100000111110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100000111110011) && ({row_reg, col_reg}<16'b0100000111110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000111110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000111110111) && ({row_reg, col_reg}<16'b0100000111111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100000111111110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}==16'b0100000111111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100001000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001000000001) && ({row_reg, col_reg}<16'b0100001000000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100001000000100) && ({row_reg, col_reg}<16'b0100001000001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001000001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100001000001001) && ({row_reg, col_reg}<16'b0100001000001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001000001100) && ({row_reg, col_reg}<16'b0100001000001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001000001110) && ({row_reg, col_reg}<16'b0100001000010001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100001000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100001000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001000010011) && ({row_reg, col_reg}<16'b0100001000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100001000100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001000100110) && ({row_reg, col_reg}<16'b0100001000101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001000101001) && ({row_reg, col_reg}<16'b0100001000101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001000101011) && ({row_reg, col_reg}<16'b0100001000101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100001000101101) && ({row_reg, col_reg}<16'b0100001000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001000110000) && ({row_reg, col_reg}<16'b0100001000110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100001000110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001000110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001000110100) && ({row_reg, col_reg}<16'b0100001000110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100001000110111) && ({row_reg, col_reg}<16'b0100001000111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100001000111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100001000111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001000111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100001000111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100001000111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100001000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001000111111) && ({row_reg, col_reg}<16'b0100001001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001001000001) && ({row_reg, col_reg}<16'b0100001001000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100001001000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001001000100) && ({row_reg, col_reg}<16'b0100001001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001001000111) && ({row_reg, col_reg}<16'b0100001001001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001001001010) && ({row_reg, col_reg}<16'b0100001001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001001001100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0100001001001101) && ({row_reg, col_reg}<16'b0100001001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001001001111) && ({row_reg, col_reg}<16'b0100001001010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100001001010011) && ({row_reg, col_reg}<16'b0100001001010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100001001010110) && ({row_reg, col_reg}<16'b0100001001011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100001001011001) && ({row_reg, col_reg}<16'b0100001001011011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100001001011011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100001001011100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0100001001011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100001001011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001001011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001001100000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0100001001100001) && ({row_reg, col_reg}<16'b0100001001100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100001001100011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0100001001100100) && ({row_reg, col_reg}<16'b0100001001100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001001100111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100001001101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100001001101001) && ({row_reg, col_reg}<16'b0100001001101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100001001101101) && ({row_reg, col_reg}<16'b0100001001110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001001110001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0100001001110010) && ({row_reg, col_reg}<16'b0100001001110100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0100001001110100) && ({row_reg, col_reg}<16'b0100001001110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001001110110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100001001110111) && ({row_reg, col_reg}<16'b0100001001111001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100001001111001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0100001001111010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0100001001111011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0100001001111100) && ({row_reg, col_reg}<16'b0100001001111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001001111110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100001001111111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100001010000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100001010000001) && ({row_reg, col_reg}<16'b0100001010000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100001010000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100001010000100) && ({row_reg, col_reg}<16'b0100001010000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100001010000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001010000111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0100001010001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100001010001001) && ({row_reg, col_reg}<16'b0100001010001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001010001011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100001010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001010001101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100001010001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001010001111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100001010010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001010010001)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0100001010010010) && ({row_reg, col_reg}<16'b0100001010010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001010010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100001010010111) && ({row_reg, col_reg}<16'b0100001010011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100001010011001) && ({row_reg, col_reg}<16'b0100001010011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001010011011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100001010011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100001010011101) && ({row_reg, col_reg}<16'b0100001010100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001010100000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100001010100001) && ({row_reg, col_reg}<16'b0100001010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100001010100011) && ({row_reg, col_reg}<16'b0100001010100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100001010100111) && ({row_reg, col_reg}<16'b0100001010101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100001010101011) && ({row_reg, col_reg}<16'b0100001010101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100001010101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100001010101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001010101111) && ({row_reg, col_reg}<16'b0100001010110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001010110001)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0100001010110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100001010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001010110101) && ({row_reg, col_reg}<16'b0100001010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001010111101) && ({row_reg, col_reg}<16'b0100001011000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100001011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100001011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001011000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100001011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100001011000100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100001011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100001011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001011000111) && ({row_reg, col_reg}<16'b0100001011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001011001111) && ({row_reg, col_reg}<16'b0100001011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001011010001) && ({row_reg, col_reg}<16'b0100001011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100001011110000) && ({row_reg, col_reg}<16'b0100001011110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001011110010) && ({row_reg, col_reg}<16'b0100001011110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001011110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001011110111) && ({row_reg, col_reg}<16'b0100001011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100001011111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001011111011) && ({row_reg, col_reg}<16'b0100001011111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100001011111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100001011111110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}==16'b0100001011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001100000000) && ({row_reg, col_reg}<16'b0100001100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001100000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100001100000111) && ({row_reg, col_reg}<16'b0100001100001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001100001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100001100001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100001100001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100001100001100) && ({row_reg, col_reg}<16'b0100001100001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001100001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001100001111) && ({row_reg, col_reg}<16'b0100001100010001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100001100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100001100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001100010011) && ({row_reg, col_reg}<16'b0100001100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100001100100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001100100110) && ({row_reg, col_reg}<16'b0100001100101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100001100101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001100101011) && ({row_reg, col_reg}<16'b0100001100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100001100101101) && ({row_reg, col_reg}<16'b0100001100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001100110000) && ({row_reg, col_reg}<16'b0100001100110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001100110010) && ({row_reg, col_reg}<16'b0100001100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001100110100) && ({row_reg, col_reg}<16'b0100001100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100001100110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100001100110111) && ({row_reg, col_reg}<16'b0100001100111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001100111001) && ({row_reg, col_reg}<16'b0100001100111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100001100111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001100111101) && ({row_reg, col_reg}<16'b0100001100111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100001100111111) && ({row_reg, col_reg}<16'b0100001101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001101000001) && ({row_reg, col_reg}<16'b0100001101000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100001101000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001101000100) && ({row_reg, col_reg}<16'b0100001101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001101000111) && ({row_reg, col_reg}<16'b0100001101001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100001101001001) && ({row_reg, col_reg}<16'b0100001101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100001101001100) && ({row_reg, col_reg}<16'b0100001101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001101001111) && ({row_reg, col_reg}<16'b0100001101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001101010100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100001101010101) && ({row_reg, col_reg}<16'b0100001101010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100001101010111) && ({row_reg, col_reg}<16'b0100001101011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001101011001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100001101011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100001101011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001101011100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0100001101011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100001101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001101011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0100001101100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100001101100001) && ({row_reg, col_reg}<16'b0100001101100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100001101100011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0100001101100100) && ({row_reg, col_reg}<16'b0100001101100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001101100110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100001101100111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100001101101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001101101001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100001101101010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100001101101011) && ({row_reg, col_reg}<16'b0100001101101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100001101101101) && ({row_reg, col_reg}<16'b0100001101110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100001101110010) && ({row_reg, col_reg}<16'b0100001101110100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0100001101110100) && ({row_reg, col_reg}<16'b0100001101110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001101110110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100001101110111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0100001101111000) && ({row_reg, col_reg}<16'b0100001101111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100001101111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100001101111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001101111101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100001101111110) && ({row_reg, col_reg}<16'b0100001110000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100001110000000)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0100001110000001)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0100001110000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001110000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100001110000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001110000101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100001110000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001110000111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0100001110001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001110001001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100001110001010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001110001011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0100001110001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001110001101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100001110001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001110001111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100001110010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001110010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100001110010010) && ({row_reg, col_reg}<16'b0100001110010100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0100001110010100) && ({row_reg, col_reg}<16'b0100001110010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001110010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100001110010111) && ({row_reg, col_reg}<16'b0100001110011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001110011001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100001110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001110011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100001110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100001110011101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0100001110011110) && ({row_reg, col_reg}<16'b0100001110100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001110100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001110100001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0100001110100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001110100011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100001110100100) && ({row_reg, col_reg}<16'b0100001110100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100001110100111) && ({row_reg, col_reg}<16'b0100001110101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100001110101001) && ({row_reg, col_reg}<16'b0100001110101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001110101011) && ({row_reg, col_reg}<16'b0100001110101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100001110101101) && ({row_reg, col_reg}<16'b0100001110101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001110101111) && ({row_reg, col_reg}<16'b0100001110110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001110110101) && ({row_reg, col_reg}<16'b0100001110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001110111101) && ({row_reg, col_reg}<16'b0100001110111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001110111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001111000000) && ({row_reg, col_reg}<16'b0100001111000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001111000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100001111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100001111000100) && ({row_reg, col_reg}<16'b0100001111000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001111000111) && ({row_reg, col_reg}<16'b0100001111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001111001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001111001111) && ({row_reg, col_reg}<16'b0100001111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001111010001) && ({row_reg, col_reg}<16'b0100001111110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100001111110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001111110001) && ({row_reg, col_reg}<16'b0100001111111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001111111011) && ({row_reg, col_reg}<16'b0100001111111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0100001111111110) && ({row_reg, col_reg}<16'b0100010000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010000000000) && ({row_reg, col_reg}<16'b0100010000000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010000000011) && ({row_reg, col_reg}<16'b0100010000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010000000101) && ({row_reg, col_reg}<16'b0100010000000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100010000000111) && ({row_reg, col_reg}<16'b0100010000001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010000001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100010000001011) && ({row_reg, col_reg}<16'b0100010000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010000001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100010000010000) && ({row_reg, col_reg}<16'b0100010000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010000010011) && ({row_reg, col_reg}<16'b0100010000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010000100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010000100110) && ({row_reg, col_reg}<16'b0100010000101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010000101000) && ({row_reg, col_reg}<16'b0100010000101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010000101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010000101011) && ({row_reg, col_reg}<16'b0100010000101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010000101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100010000101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010000101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010000110000) && ({row_reg, col_reg}<16'b0100010000110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010000110010) && ({row_reg, col_reg}<16'b0100010000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010000110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100010000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100010000110111) && ({row_reg, col_reg}<16'b0100010000111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010000111001) && ({row_reg, col_reg}<16'b0100010000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100010000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010000111111) && ({row_reg, col_reg}<16'b0100010001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100010001000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100010001000010) && ({row_reg, col_reg}<16'b0100010001000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010001000100) && ({row_reg, col_reg}<16'b0100010001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010001000111) && ({row_reg, col_reg}<16'b0100010001001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100010001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100010001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010001001100) && ({row_reg, col_reg}<16'b0100010001001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100010001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100010001001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010001010000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0100010001010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100010001010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100010001010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100010001010100) && ({row_reg, col_reg}<16'b0100010001010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100010001010111) && ({row_reg, col_reg}<16'b0100010001011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010001011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100010001011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100010001011011) && ({row_reg, col_reg}<16'b0100010001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100010001011111) && ({row_reg, col_reg}<16'b0100010001100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100010001100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100010001100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100010001100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100010001100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100010001100101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100010001100110) && ({row_reg, col_reg}<16'b0100010001101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100010001101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010001101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010001101011) && ({row_reg, col_reg}<16'b0100010001101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100010001101101) && ({row_reg, col_reg}<16'b0100010001110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100010001110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100010001110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100010001110010) && ({row_reg, col_reg}<16'b0100010001110110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0100010001110110) && ({row_reg, col_reg}<16'b0100010001111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100010001111000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0100010001111001) && ({row_reg, col_reg}<16'b0100010001111100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0100010001111100) && ({row_reg, col_reg}<16'b0100010001111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100010001111111)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0100010010000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100010010000001) && ({row_reg, col_reg}<16'b0100010010000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010010000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100010010000101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100010010000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100010010000111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0100010010001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010010001001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100010010001010) && ({row_reg, col_reg}<16'b0100010010001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100010010001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100010010001110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0100010010001111) && ({row_reg, col_reg}<16'b0100010010010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010010010001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0100010010010010) && ({row_reg, col_reg}<16'b0100010010010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100010010010101) && ({row_reg, col_reg}<16'b0100010010010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100010010010111) && ({row_reg, col_reg}<16'b0100010010011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100010010011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100010010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100010010011101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0100010010011110) && ({row_reg, col_reg}<16'b0100010010100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010010100000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0100010010100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100010010100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010010100011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100010010100100) && ({row_reg, col_reg}<16'b0100010010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100010010100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0100010010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100010010101000) && ({row_reg, col_reg}<16'b0100010010101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010010101010) && ({row_reg, col_reg}<16'b0100010010110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010010110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100010010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100010010110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010010110111) && ({row_reg, col_reg}<16'b0100010010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010010111101) && ({row_reg, col_reg}<16'b0100010010111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010010111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100010011000000) && ({row_reg, col_reg}<16'b0100010011000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010011000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100010011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100010011000100) && ({row_reg, col_reg}<16'b0100010011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010011000110) && ({row_reg, col_reg}<16'b0100010011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100010011001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010011010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010011010001) && ({row_reg, col_reg}<16'b0100010011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100010011110000) && ({row_reg, col_reg}<16'b0100010011110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010011110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100010011110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010011110111) && ({row_reg, col_reg}<16'b0100010011111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100010011111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010011111011) && ({row_reg, col_reg}<16'b0100010011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010011111110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}==16'b0100010011111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010100000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010100000001) && ({row_reg, col_reg}<16'b0100010100000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010100000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010100000100) && ({row_reg, col_reg}<16'b0100010100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010100010011) && ({row_reg, col_reg}<16'b0100010100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010100100100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100010100100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010100100110) && ({row_reg, col_reg}<16'b0100010100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010100101000) && ({row_reg, col_reg}<16'b0100010100101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010100101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010100101011) && ({row_reg, col_reg}<16'b0100010100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010100101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100010100101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010100101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100010100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010100110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010100110010) && ({row_reg, col_reg}<16'b0100010100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010100110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100010100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010100110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100010100110111) && ({row_reg, col_reg}<16'b0100010100111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100010100111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100010100111010) && ({row_reg, col_reg}<16'b0100010100111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010100111100) && ({row_reg, col_reg}<16'b0100010100111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100010100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010100111111) && ({row_reg, col_reg}<16'b0100010101000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100010101000010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100010101000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010101000100) && ({row_reg, col_reg}<16'b0100010101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010101000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100010101000111) && ({row_reg, col_reg}<16'b0100010101001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100010101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100010101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010101001100) && ({row_reg, col_reg}<16'b0100010101001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100010101001110) && ({row_reg, col_reg}<16'b0100010101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100010101010000) && ({row_reg, col_reg}<16'b0100010101010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100010101010010) && ({row_reg, col_reg}<16'b0100010101010100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0100010101010100) && ({row_reg, col_reg}<16'b0100010101010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100010101010111) && ({row_reg, col_reg}<16'b0100010101011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100010101011001) && ({row_reg, col_reg}<16'b0100010101011011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100010101011011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0100010101011100) && ({row_reg, col_reg}<16'b0100010101011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010101011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0100010101100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100010101100001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0100010101100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100010101100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100010101100100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100010101100101) && ({row_reg, col_reg}<16'b0100010101100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010101100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100010101101000) && ({row_reg, col_reg}<16'b0100010101101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010101101011) && ({row_reg, col_reg}<16'b0100010101101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100010101101101) && ({row_reg, col_reg}<16'b0100010101101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100010101101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010101110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100010101110001) && ({row_reg, col_reg}<16'b0100010101110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100010101110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0100010101110110) && ({row_reg, col_reg}<16'b0100010101111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100010101111000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100010101111001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0100010101111010) && ({row_reg, col_reg}<16'b0100010101111100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100010101111100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100010101111101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100010101111110)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0100010101111111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100010110000000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0100010110000001) && ({row_reg, col_reg}<16'b0100010110000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010110000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100010110000101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0100010110000110) && ({row_reg, col_reg}<16'b0100010110001000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100010110001000) && ({row_reg, col_reg}<16'b0100010110001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010110001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100010110001101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100010110001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100010110001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010110010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100010110010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010110010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100010110010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100010110010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100010110010101) && ({row_reg, col_reg}<16'b0100010110010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100010110010111) && ({row_reg, col_reg}<16'b0100010110011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100010110011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100010110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100010110011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100010110011110) && ({row_reg, col_reg}<16'b0100010110100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100010110100011) && ({row_reg, col_reg}<16'b0100010110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100010110100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0100010110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010110101000) && ({row_reg, col_reg}<16'b0100010110101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100010110101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010110101011) && ({row_reg, col_reg}<16'b0100010110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010110110100) && ({row_reg, col_reg}<16'b0100010110110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100010110110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100010110110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010110111000) && ({row_reg, col_reg}<16'b0100010110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010110111101) && ({row_reg, col_reg}<16'b0100010110111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010110111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100010111000000) && ({row_reg, col_reg}<16'b0100010111000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010111000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100010111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010111000100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010111000101) && ({row_reg, col_reg}<16'b0100010111001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010111001010) && ({row_reg, col_reg}<16'b0100010111001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100010111001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010111010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010111010001) && ({row_reg, col_reg}<16'b0100010111110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100010111110000) && ({row_reg, col_reg}<16'b0100010111110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010111110100) && ({row_reg, col_reg}<16'b0100010111110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010111110110) && ({row_reg, col_reg}<16'b0100010111111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100010111111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010111111011) && ({row_reg, col_reg}<16'b0100010111111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010111111110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0100010111111111) && ({row_reg, col_reg}<16'b0100011000000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011000000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100011000000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100011000000011) && ({row_reg, col_reg}<16'b0100011000000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011000000110) && ({row_reg, col_reg}<16'b0100011000001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011000001001) && ({row_reg, col_reg}<16'b0100011000001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011000001100) && ({row_reg, col_reg}<16'b0100011000001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011000001110) && ({row_reg, col_reg}<16'b0100011000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011000010011) && ({row_reg, col_reg}<16'b0100011000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100011000100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011000100110) && ({row_reg, col_reg}<16'b0100011000101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011000101000) && ({row_reg, col_reg}<16'b0100011000101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011000101011) && ({row_reg, col_reg}<16'b0100011000101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011000101101) && ({row_reg, col_reg}<16'b0100011000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011000110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011000110010) && ({row_reg, col_reg}<16'b0100011000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011000110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100011000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011000110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100011000110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100011000111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100011000111001) && ({row_reg, col_reg}<16'b0100011000111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100011000111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011000111100) && ({row_reg, col_reg}<16'b0100011000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100011000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011000111111) && ({row_reg, col_reg}<16'b0100011001000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100011001000010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100011001000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011001000100) && ({row_reg, col_reg}<16'b0100011001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011001000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100011001000111) && ({row_reg, col_reg}<16'b0100011001001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100011001001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100011001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011001001100) && ({row_reg, col_reg}<16'b0100011001001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100011001001110) && ({row_reg, col_reg}<16'b0100011001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100011001010000) && ({row_reg, col_reg}<16'b0100011001010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100011001010011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0100011001010100) && ({row_reg, col_reg}<16'b0100011001010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011001010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100011001011000) && ({row_reg, col_reg}<16'b0100011001011011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011001011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100011001011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100011001011101) && ({row_reg, col_reg}<16'b0100011001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011001011111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100011001100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100011001100001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0100011001100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100011001100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100011001100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100011001100101) && ({row_reg, col_reg}<16'b0100011001100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100011001100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100011001101000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100011001101001) && ({row_reg, col_reg}<16'b0100011001101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100011001101011) && ({row_reg, col_reg}<16'b0100011001101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100011001101101) && ({row_reg, col_reg}<16'b0100011001101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100011001101111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100011001110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100011001110001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100011001110010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0100011001110011) && ({row_reg, col_reg}<16'b0100011001110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100011001110101) && ({row_reg, col_reg}<16'b0100011001111001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0100011001111001) && ({row_reg, col_reg}<16'b0100011001111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100011001111011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100011001111100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0100011001111101) && ({row_reg, col_reg}<16'b0100011010000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100011010000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100011010000001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100011010000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011010000011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100011010000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100011010000101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100011010000110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100011010000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100011010001000) && ({row_reg, col_reg}<16'b0100011010001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100011010001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100011010001110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100011010001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011010010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100011010010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011010010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100011010010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100011010010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100011010010101) && ({row_reg, col_reg}<16'b0100011010010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011010010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011010011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100011010011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100011010011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100011010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100011010011101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100011010011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011010011111) && ({row_reg, col_reg}<16'b0100011010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100011010100011) && ({row_reg, col_reg}<16'b0100011010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011010100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0100011010100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011010101000) && ({row_reg, col_reg}<16'b0100011010101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100011010101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011010101011) && ({row_reg, col_reg}<16'b0100011010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011010110100) && ({row_reg, col_reg}<16'b0100011010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011010110110) && ({row_reg, col_reg}<16'b0100011010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100011010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011010111001) && ({row_reg, col_reg}<16'b0100011010111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011010111110) && ({row_reg, col_reg}<16'b0100011011000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100011011000000) && ({row_reg, col_reg}<16'b0100011011000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011011000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100011011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100011011000100) && ({row_reg, col_reg}<16'b0100011011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011011000110) && ({row_reg, col_reg}<16'b0100011011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011011001000) && ({row_reg, col_reg}<16'b0100011011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011011001011) && ({row_reg, col_reg}<16'b0100011011001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011011001111) && ({row_reg, col_reg}<16'b0100011011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011011010001) && ({row_reg, col_reg}<16'b0100011011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100011011110000) && ({row_reg, col_reg}<16'b0100011011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011011110010) && ({row_reg, col_reg}<16'b0100011011111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100011011111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011011111011) && ({row_reg, col_reg}<16'b0100011011111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0100011011111110) && ({row_reg, col_reg}<16'b0100011100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011100000000) && ({row_reg, col_reg}<16'b0100011100000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011100000100) && ({row_reg, col_reg}<16'b0100011100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011100000111) && ({row_reg, col_reg}<16'b0100011100001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011100001001) && ({row_reg, col_reg}<16'b0100011100001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011100001100) && ({row_reg, col_reg}<16'b0100011100001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100011100001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011100001111) && ({row_reg, col_reg}<16'b0100011100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011100010010) && ({row_reg, col_reg}<16'b0100011100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100011100100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011100100110) && ({row_reg, col_reg}<16'b0100011100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011100101000) && ({row_reg, col_reg}<16'b0100011100101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011100101010) && ({row_reg, col_reg}<16'b0100011100101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011100101101) && ({row_reg, col_reg}<16'b0100011100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011100110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100011100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100011100110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100011100111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100011100111001) && ({row_reg, col_reg}<16'b0100011100111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011100111100) && ({row_reg, col_reg}<16'b0100011100111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100011100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011100111111) && ({row_reg, col_reg}<16'b0100011101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100011101000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100011101000100) && ({row_reg, col_reg}<16'b0100011101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011101000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100011101000111) && ({row_reg, col_reg}<16'b0100011101001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100011101001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100011101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100011101001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100011101001101) && ({row_reg, col_reg}<16'b0100011101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011101001111) && ({row_reg, col_reg}<16'b0100011101010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011101010101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100011101010110) && ({row_reg, col_reg}<16'b0100011101011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100011101011000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100011101011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011101011010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0100011101011011) && ({row_reg, col_reg}<16'b0100011101011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100011101011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011101011110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0100011101011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011101100000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100011101100001)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0100011101100010) && ({row_reg, col_reg}<16'b0100011101100100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100011101100100)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0100011101100101)) color_data = 12'b100001110101;
		if(({row_reg, col_reg}==16'b0100011101100110)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0100011101100111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100011101101000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100011101101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100011101101010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0100011101101011) && ({row_reg, col_reg}<16'b0100011101101101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100011101101101) && ({row_reg, col_reg}<16'b0100011101101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100011101101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100011101110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100011101110001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100011101110010)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}>=16'b0100011101110011) && ({row_reg, col_reg}<16'b0100011101110101)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==16'b0100011101110101)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0100011101110110)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0100011101110111) && ({row_reg, col_reg}<16'b0100011101111001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100011101111001) && ({row_reg, col_reg}<16'b0100011101111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100011101111011)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0100011101111100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100011101111101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100011101111110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0100011101111111)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0100011110000000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0100011110000001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0100011110000010) && ({row_reg, col_reg}<16'b0100011110000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100011110000100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0100011110000101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100011110000110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100011110000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100011110001000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011110001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100011110001010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100011110001011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100011110001100)) color_data = 12'b100001110101;
		if(({row_reg, col_reg}==16'b0100011110001101)) color_data = 12'b100110000110;
		if(({row_reg, col_reg}==16'b0100011110001110)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==16'b0100011110001111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100011110010000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100011110010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100011110010010) && ({row_reg, col_reg}<16'b0100011110010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011110010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011110011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100011110011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100011110011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100011110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100011110011101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100011110011110) && ({row_reg, col_reg}<16'b0100011110100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011110100000) && ({row_reg, col_reg}<16'b0100011110100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100011110100011) && ({row_reg, col_reg}<16'b0100011110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011110100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0100011110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100011110101000) && ({row_reg, col_reg}<16'b0100011110101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011110101011) && ({row_reg, col_reg}<16'b0100011110110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100011110110000) && ({row_reg, col_reg}<16'b0100011110110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100011110110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011110110100) && ({row_reg, col_reg}<16'b0100011110110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011110110110) && ({row_reg, col_reg}<16'b0100011110111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100011110111001) && ({row_reg, col_reg}<16'b0100011110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011110111101) && ({row_reg, col_reg}<16'b0100011110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100011110111111) && ({row_reg, col_reg}<16'b0100011111000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100011111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011111000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100011111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100011111000100) && ({row_reg, col_reg}<16'b0100011111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011111000110) && ({row_reg, col_reg}<16'b0100011111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011111001000) && ({row_reg, col_reg}<16'b0100011111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011111001011) && ({row_reg, col_reg}<16'b0100011111001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011111001111) && ({row_reg, col_reg}<16'b0100011111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011111010001) && ({row_reg, col_reg}<16'b0100011111110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100011111110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011111110001) && ({row_reg, col_reg}<16'b0100011111110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100011111110011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=16'b0100011111110100) && ({row_reg, col_reg}<16'b0100011111110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100011111110110) && ({row_reg, col_reg}<16'b0100011111111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100011111111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100011111111001) && ({row_reg, col_reg}<16'b0100011111111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011111111011) && ({row_reg, col_reg}<16'b0100011111111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0100011111111110) && ({row_reg, col_reg}<16'b0100100000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100000000000) && ({row_reg, col_reg}<16'b0100100000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100000000110) && ({row_reg, col_reg}<16'b0100100000001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100000001000) && ({row_reg, col_reg}<16'b0100100000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100000001101) && ({row_reg, col_reg}<16'b0100100000001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100000001111) && ({row_reg, col_reg}<16'b0100100000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100100000010010) && ({row_reg, col_reg}<16'b0100100000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100100000100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100000100110) && ({row_reg, col_reg}<16'b0100100000101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100000101000) && ({row_reg, col_reg}<16'b0100100000101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100000101010) && ({row_reg, col_reg}<16'b0100100000101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100100000101101) && ({row_reg, col_reg}<16'b0100100000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100000110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100100000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100100000110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100100000111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100100000111001) && ({row_reg, col_reg}<16'b0100100000111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100000111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100000111100) && ({row_reg, col_reg}<16'b0100100000111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100100000111111) && ({row_reg, col_reg}<16'b0100100001000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100001000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100100001000100) && ({row_reg, col_reg}<16'b0100100001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100100001000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100100001000111) && ({row_reg, col_reg}<16'b0100100001001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100001001010) && ({row_reg, col_reg}<16'b0100100001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100100001001100) && ({row_reg, col_reg}<16'b0100100001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100001001111) && ({row_reg, col_reg}<16'b0100100001010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100100001010101) && ({row_reg, col_reg}<16'b0100100001011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100001011001) && ({row_reg, col_reg}<16'b0100100001011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100100001011011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0100100001011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100100001011101) && ({row_reg, col_reg}<16'b0100100001011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100100001011111) && ({row_reg, col_reg}<16'b0100100001100001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100100001100001)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100100001100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100100001100011)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0100100001100100)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}>=16'b0100100001100101) && ({row_reg, col_reg}<16'b0100100001100111)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0100100001100111)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0100100001101000)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}>=16'b0100100001101001) && ({row_reg, col_reg}<16'b0100100001101100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100100001101100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100100001101101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100100001101110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100100001101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100100001110000)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0100100001110001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0100100001110010)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0100100001110011)) color_data = 12'b101111001001;
		if(({row_reg, col_reg}==16'b0100100001110100)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0100100001110101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0100100001110110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100100001110111) && ({row_reg, col_reg}<16'b0100100001111100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100100001111100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100100001111101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0100100001111110)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0100100001111111)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0100100010000000)) color_data = 12'b101010111001;
		if(({row_reg, col_reg}==16'b0100100010000001)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0100100010000010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=16'b0100100010000011) && ({row_reg, col_reg}<16'b0100100010000101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100100010000101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100100010000110)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100100010000111)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0100100010001000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100100010001001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100100010001010)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0100100010001011)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0100100010001100)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0100100010001101)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0100100010001110)) color_data = 12'b100110101000;
		if(({row_reg, col_reg}==16'b0100100010001111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0100100010010000)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0100100010010001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100100010010010)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0100100010010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100100010010100) && ({row_reg, col_reg}<16'b0100100010010110)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0100100010010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100010010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100010011000) && ({row_reg, col_reg}<16'b0100100010011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100100010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100100010011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100100010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100100010011101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100100010011110) && ({row_reg, col_reg}<16'b0100100010100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100010100000) && ({row_reg, col_reg}<16'b0100100010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100100010100011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100100010100100) && ({row_reg, col_reg}<16'b0100100010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100100010100110) && ({row_reg, col_reg}<16'b0100100010110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100100010110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100010110001) && ({row_reg, col_reg}<16'b0100100010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100100010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100100010110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100100010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100010110110) && ({row_reg, col_reg}<16'b0100100010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100100010111000) && ({row_reg, col_reg}<16'b0100100010111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100100010111010) && ({row_reg, col_reg}<16'b0100100010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100010111100)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==16'b0100100010111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100100010111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100100010111111) && ({row_reg, col_reg}<16'b0100100011000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100100011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100011000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100100011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100100011000100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100100011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100100011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100100011000111) && ({row_reg, col_reg}<16'b0100100011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100011001001) && ({row_reg, col_reg}<16'b0100100011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100011001011) && ({row_reg, col_reg}<16'b0100100011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100100011001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100100011001111) && ({row_reg, col_reg}<16'b0100100011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100011010001) && ({row_reg, col_reg}<16'b0100100011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100100011110000) && ({row_reg, col_reg}<16'b0100100011110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100011110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100011110100) && ({row_reg, col_reg}<16'b0100100011111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100100011111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100011111011) && ({row_reg, col_reg}<16'b0100100011111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0100100011111110) && ({row_reg, col_reg}<16'b0100100100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100100000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100100100000001) && ({row_reg, col_reg}<16'b0100100100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100100000110) && ({row_reg, col_reg}<16'b0100100100001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100100001000) && ({row_reg, col_reg}<16'b0100100100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100100001110) && ({row_reg, col_reg}<16'b0100100100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100100010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100100100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100100010010) && ({row_reg, col_reg}<16'b0100100100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100100100100100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100100100100101) && ({row_reg, col_reg}<16'b0100100100100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100100100111) && ({row_reg, col_reg}<16'b0100100100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100100101001) && ({row_reg, col_reg}<16'b0100100100101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100100100101011) && ({row_reg, col_reg}<16'b0100100100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100100100101101) && ({row_reg, col_reg}<16'b0100100100110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100100110010) && ({row_reg, col_reg}<16'b0100100100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100100110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100100100110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100100100111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100100100111001) && ({row_reg, col_reg}<16'b0100100100111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100100111100) && ({row_reg, col_reg}<16'b0100100100111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100100100111111) && ({row_reg, col_reg}<16'b0100100101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100101000100) && ({row_reg, col_reg}<16'b0100100101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100100101000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100100101000111) && ({row_reg, col_reg}<16'b0100100101001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100101001010) && ({row_reg, col_reg}<16'b0100100101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100100101001100) && ({row_reg, col_reg}<16'b0100100101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100101001111) && ({row_reg, col_reg}<16'b0100100101011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100100101011000) && ({row_reg, col_reg}<16'b0100100101011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100101011010) && ({row_reg, col_reg}<16'b0100100101011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100100101011100) && ({row_reg, col_reg}<16'b0100100101011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100100101011111) && ({row_reg, col_reg}<16'b0100100101100010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100100101100010)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100100101100011)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0100100101100100)) color_data = 12'b100110101000;
		if(({row_reg, col_reg}==16'b0100100101100101)) color_data = 12'b101111001001;
		if(({row_reg, col_reg}==16'b0100100101100110)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==16'b0100100101100111)) color_data = 12'b101010111000;
		if(({row_reg, col_reg}==16'b0100100101101000)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0100100101101001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0100100101101010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=16'b0100100101101011) && ({row_reg, col_reg}<16'b0100100101101101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100100101101101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100100101101110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100100101101111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100100101110000)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0100100101110001)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0100100101110010)) color_data = 12'b101111001001;
		if(({row_reg, col_reg}==16'b0100100101110011)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==16'b0100100101110100)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0100100101110101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100100101110110)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100100101110111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100100101111000)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100100101111001) && ({row_reg, col_reg}<16'b0100100101111011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100100101111011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100100101111100)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0100100101111101)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=16'b0100100101111110) && ({row_reg, col_reg}<16'b0100100110000000)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==16'b0100100110000000)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0100100110000001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0100100110000010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0100100110000011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100100110000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100100110000101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100100110000110)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100100110000111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100100110001000)) color_data = 12'b011110000110;
		if(({row_reg, col_reg}>=16'b0100100110001001) && ({row_reg, col_reg}<16'b0100100110001011)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0100100110001011)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}>=16'b0100100110001100) && ({row_reg, col_reg}<16'b0100100110001110)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==16'b0100100110001110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0100100110001111)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100100110010000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0100100110010001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100100110010010)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0100100110010011)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0100100110010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100110010101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0100100110010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100100110010111) && ({row_reg, col_reg}<16'b0100100110011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100100110011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100100110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100100110011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100100110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100100110011101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100100110011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100100110011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100110100000) && ({row_reg, col_reg}<16'b0100100110100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100100110100011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100100110100100) && ({row_reg, col_reg}<16'b0100100110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100100110100110) && ({row_reg, col_reg}<16'b0100100110110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100100110110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100100110110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100100110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100110110100) && ({row_reg, col_reg}<16'b0100100110110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100100110110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100100110110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100100110111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100100110111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100100110111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100110111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100110111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100100110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100100110111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100100110111111) && ({row_reg, col_reg}<16'b0100100111000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100111000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100100111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100100111000100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100100111000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100100111000110) && ({row_reg, col_reg}<16'b0100100111001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100100111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100111001001) && ({row_reg, col_reg}<16'b0100100111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100111001011) && ({row_reg, col_reg}<16'b0100100111001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100100111001101) && ({row_reg, col_reg}<16'b0100100111001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100100111001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100100111010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100111010001) && ({row_reg, col_reg}<16'b0100100111110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100100111110000) && ({row_reg, col_reg}<16'b0100100111110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100111110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100111110100) && ({row_reg, col_reg}<16'b0100100111111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100100111111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100111111011) && ({row_reg, col_reg}<16'b0100100111111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0100100111111110) && ({row_reg, col_reg}<16'b0100101000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101000000000) && ({row_reg, col_reg}<16'b0100101000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101000000110) && ({row_reg, col_reg}<16'b0100101000001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101000001001) && ({row_reg, col_reg}<16'b0100101000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101000010011) && ({row_reg, col_reg}<16'b0100101000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100101000100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100101000100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101000100111) && ({row_reg, col_reg}<16'b0100101000101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100101000101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101000101010) && ({row_reg, col_reg}<16'b0100101000101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101000101110) && ({row_reg, col_reg}<16'b0100101000110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101000110010) && ({row_reg, col_reg}<16'b0100101000110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100101000110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100101000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101000110110) && ({row_reg, col_reg}<16'b0100101000111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101000111001) && ({row_reg, col_reg}<16'b0100101000111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100101000111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101000111100) && ({row_reg, col_reg}<16'b0100101000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100101000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101000111111) && ({row_reg, col_reg}<16'b0100101001000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101001000100) && ({row_reg, col_reg}<16'b0100101001000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101001000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100101001001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100101001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101001001010) && ({row_reg, col_reg}<16'b0100101001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100101001001100) && ({row_reg, col_reg}<16'b0100101001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101001001111) && ({row_reg, col_reg}<16'b0100101001011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100101001011000) && ({row_reg, col_reg}<16'b0100101001011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101001011010) && ({row_reg, col_reg}<16'b0100101001011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101001011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100101001011110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100101001011111)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0100101001100000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100101001100001) && ({row_reg, col_reg}<16'b0100101001100011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100101001100011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100101001100100)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0100101001100101)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==16'b0100101001100110)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0100101001100111)) color_data = 12'b110011001001;
		if(({row_reg, col_reg}==16'b0100101001101000)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0100101001101001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=16'b0100101001101010) && ({row_reg, col_reg}<16'b0100101001101101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100101001101101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100101001101110)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100101001101111)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0100101001110000)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0100101001110001)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0100101001110010)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==16'b0100101001110011)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0100101001110100)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0100101001110101)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}>=16'b0100101001110110) && ({row_reg, col_reg}<16'b0100101001111010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100101001111010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100101001111011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0100101001111100)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==16'b0100101001111101)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0100101001111110)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0100101001111111)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0100101010000000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0100101010000001)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0100101010000010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0100101010000011) && ({row_reg, col_reg}<16'b0100101010000110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100101010000110)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0100101010000111)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==16'b0100101010001000)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0100101010001001)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0100101010001010)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0100101010001011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=16'b0100101010001100) && ({row_reg, col_reg}<16'b0100101010001110)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}>=16'b0100101010001110) && ({row_reg, col_reg}<16'b0100101010010000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100101010010000)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0100101010010001)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0100101010010010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100101010010011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100101010010100) && ({row_reg, col_reg}<16'b0100101010010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100101010010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100101010011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101010011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100101010011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100101010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100101010011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100101010011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101010011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100101010100000) && ({row_reg, col_reg}<16'b0100101010100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100101010100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101010100011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100101010100100) && ({row_reg, col_reg}<16'b0100101010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100101010100110) && ({row_reg, col_reg}<16'b0100101010101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101010101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100101010101010) && ({row_reg, col_reg}<16'b0100101010101101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100101010101101) && ({row_reg, col_reg}<16'b0100101010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101010110100) && ({row_reg, col_reg}<16'b0100101010110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100101010110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100101010110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101010111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100101010111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100101010111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101010111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101010111100) && ({row_reg, col_reg}<16'b0100101010111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100101010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101011000000) && ({row_reg, col_reg}<16'b0100101011000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101011000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100101011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101011000100) && ({row_reg, col_reg}<16'b0100101011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101011000110) && ({row_reg, col_reg}<16'b0100101011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101011001001) && ({row_reg, col_reg}<16'b0100101011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101011001011) && ({row_reg, col_reg}<16'b0100101011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100101011001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100101011001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100101011010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101011010001) && ({row_reg, col_reg}<16'b0100101011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101011110000) && ({row_reg, col_reg}<16'b0100101011110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101011110011) && ({row_reg, col_reg}<16'b0100101011110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101011110101) && ({row_reg, col_reg}<16'b0100101011111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100101011111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101011111011) && ({row_reg, col_reg}<16'b0100101011111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0100101011111110) && ({row_reg, col_reg}<16'b0100101100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101100000000) && ({row_reg, col_reg}<16'b0100101100000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101100000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101100000101) && ({row_reg, col_reg}<16'b0100101100000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101100000111) && ({row_reg, col_reg}<16'b0100101100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101100001001) && ({row_reg, col_reg}<16'b0100101100001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101100001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101100001101) && ({row_reg, col_reg}<16'b0100101100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101100010011) && ({row_reg, col_reg}<16'b0100101100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100101100100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101100100110) && ({row_reg, col_reg}<16'b0100101100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100101100101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101100101010) && ({row_reg, col_reg}<16'b0100101100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101100101110) && ({row_reg, col_reg}<16'b0100101100110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101100110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101100110010) && ({row_reg, col_reg}<16'b0100101100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101100110100) && ({row_reg, col_reg}<16'b0100101100110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100101100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101100110111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100101100111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100101100111001) && ({row_reg, col_reg}<16'b0100101100111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100101100111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100101100111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101100111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100101100111110) && ({row_reg, col_reg}<16'b0100101101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100101101000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101101000100) && ({row_reg, col_reg}<16'b0100101101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101101000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100101101000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100101101001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100101101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101101001010) && ({row_reg, col_reg}<16'b0100101101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100101101001100) && ({row_reg, col_reg}<16'b0100101101010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101101010000) && ({row_reg, col_reg}<16'b0100101101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101101010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100101101010101) && ({row_reg, col_reg}<16'b0100101101011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100101101011000) && ({row_reg, col_reg}<16'b0100101101011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101101011010) && ({row_reg, col_reg}<16'b0100101101011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101101011101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100101101011110)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0100101101011111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0100101101100000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100101101100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0100101101100010) && ({row_reg, col_reg}<16'b0100101101100100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100101101100100)) color_data = 12'b010101100100;
		if(({row_reg, col_reg}==16'b0100101101100101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0100101101100110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==16'b0100101101100111)) color_data = 12'b101111001001;
		if(({row_reg, col_reg}==16'b0100101101101000)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0100101101101001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100101101101010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0100101101101011) && ({row_reg, col_reg}<16'b0100101101101101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100101101101101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100101101101110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100101101101111)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0100101101110000)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}>=16'b0100101101110001) && ({row_reg, col_reg}<16'b0100101101110011)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0100101101110011)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0100101101110100)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}>=16'b0100101101110101) && ({row_reg, col_reg}<16'b0100101101111001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100101101111001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100101101111010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=16'b0100101101111011) && ({row_reg, col_reg}<16'b0100101101111101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0100101101111101)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0100101101111110)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0100101101111111)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=16'b0100101110000000) && ({row_reg, col_reg}<16'b0100101110000010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100101110000010)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0100101110000011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100101110000100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0100101110000101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0100101110000110)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0100101110000111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0100101110001000)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0100101110001001)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0100101110001010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100101110001011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100101110001100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100101110001101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100101110001110)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0100101110001111)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}>=16'b0100101110010000) && ({row_reg, col_reg}<16'b0100101110010010)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0100101110010010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0100101110010011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100101110010100) && ({row_reg, col_reg}<16'b0100101110010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100101110010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101110011000) && ({row_reg, col_reg}<16'b0100101110011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100101110011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100101110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100101110011101)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0100101110011110) && ({row_reg, col_reg}<16'b0100101110100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101110100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100101110100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100101110100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101110100011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100101110100100) && ({row_reg, col_reg}<16'b0100101110100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100101110100111) && ({row_reg, col_reg}<16'b0100101110101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100101110101011) && ({row_reg, col_reg}<16'b0100101110110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100101110110000) && ({row_reg, col_reg}<16'b0100101110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101110110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100101110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101110110110) && ({row_reg, col_reg}<16'b0100101110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100101110111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100101110111001) && ({row_reg, col_reg}<16'b0100101110111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101110111011) && ({row_reg, col_reg}<16'b0100101110111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100101110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101110111110) && ({row_reg, col_reg}<16'b0100101111000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100101111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101111000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100101111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101111000100) && ({row_reg, col_reg}<16'b0100101111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101111000110) && ({row_reg, col_reg}<16'b0100101111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101111001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100101111001010)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=16'b0100101111001011) && ({row_reg, col_reg}<16'b0100101111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101111001110) && ({row_reg, col_reg}<16'b0100101111010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100101111010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101111010001) && ({row_reg, col_reg}<16'b0100101111110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101111110000) && ({row_reg, col_reg}<16'b0100101111110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101111110010) && ({row_reg, col_reg}<16'b0100101111110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101111110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100101111110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100101111110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100101111111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101111111001) && ({row_reg, col_reg}<16'b0100101111111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101111111011) && ({row_reg, col_reg}<16'b0100101111111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0100101111111110) && ({row_reg, col_reg}<16'b0100110000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100110000000000) && ({row_reg, col_reg}<16'b0100110000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110000000101) && ({row_reg, col_reg}<16'b0100110000000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110000000111) && ({row_reg, col_reg}<16'b0100110000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110000010011) && ({row_reg, col_reg}<16'b0100110000100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110000100110) && ({row_reg, col_reg}<16'b0100110000101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110000101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110000101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110000101010) && ({row_reg, col_reg}<16'b0100110000101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110000101110) && ({row_reg, col_reg}<16'b0100110000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110000110001) && ({row_reg, col_reg}<16'b0100110000110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100110000110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110000110100) && ({row_reg, col_reg}<16'b0100110000110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100110000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110000110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100110000111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100110000111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100110000111010) && ({row_reg, col_reg}<16'b0100110000111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100110000111100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0100110000111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100110000111110) && ({row_reg, col_reg}<16'b0100110001000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110001000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100110001000100) && ({row_reg, col_reg}<16'b0100110001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100110001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100110001000111) && ({row_reg, col_reg}<16'b0100110001001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110001001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100110001001010) && ({row_reg, col_reg}<16'b0100110001001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110001001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100110001001101) && ({row_reg, col_reg}<16'b0100110001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100110001001111) && ({row_reg, col_reg}<16'b0100110001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100110001010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100110001010101) && ({row_reg, col_reg}<16'b0100110001010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100110001010111) && ({row_reg, col_reg}<16'b0100110001011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110001011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100110001011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110001011101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100110001011110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0100110001011111)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0100110001100000)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==16'b0100110001100001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100110001100010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100110001100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100110001100100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100110001100101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100110001100110)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0100110001100111)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0100110001101000)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0100110001101001)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=16'b0100110001101010) && ({row_reg, col_reg}<16'b0100110001101101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100110001101101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100110001101110)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100110001101111)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0100110001110000)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0100110001110001)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0100110001110010)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0100110001110011)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0100110001110100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100110001110101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100110001110110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100110001110111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100110001111000)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0100110001111001)) color_data = 12'b011110000110;
		if(({row_reg, col_reg}==16'b0100110001111010)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0100110001111011)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0100110001111100)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0100110001111101)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0100110001111110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100110001111111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100110010000000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100110010000001) && ({row_reg, col_reg}<16'b0100110010000011)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0100110010000011)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}>=16'b0100110010000100) && ({row_reg, col_reg}<16'b0100110010000110)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==16'b0100110010000110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0100110010000111)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0100110010001000)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0100110010001001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0100110010001010) && ({row_reg, col_reg}<16'b0100110010001100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100110010001100) && ({row_reg, col_reg}<16'b0100110010001110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100110010001110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0100110010001111)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}>=16'b0100110010010000) && ({row_reg, col_reg}<16'b0100110010010010)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==16'b0100110010010010)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0100110010010011)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0100110010010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100110010010101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100110010010110) && ({row_reg, col_reg}<16'b0100110010011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100110010011000) && ({row_reg, col_reg}<16'b0100110010011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100110010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100110010011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100110010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100110010011101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0100110010011110) && ({row_reg, col_reg}<16'b0100110010100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100110010100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100110010100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100110010100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100110010100011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100110010100100) && ({row_reg, col_reg}<16'b0100110010100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100110010100111) && ({row_reg, col_reg}<16'b0100110010101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100110010101100) && ({row_reg, col_reg}<16'b0100110010110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100110010110000) && ({row_reg, col_reg}<16'b0100110010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100110010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100110010110100) && ({row_reg, col_reg}<16'b0100110010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100110010110110) && ({row_reg, col_reg}<16'b0100110010111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100110010111001) && ({row_reg, col_reg}<16'b0100110010111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100110010111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110010111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110010111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100110010111111) && ({row_reg, col_reg}<16'b0100110011000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100110011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110011000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100110011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110011000100) && ({row_reg, col_reg}<16'b0100110011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110011000110) && ({row_reg, col_reg}<16'b0100110011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110011001000) && ({row_reg, col_reg}<16'b0100110011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110011001010)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==16'b0100110011001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110011001100) && ({row_reg, col_reg}<16'b0100110011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110011001111) && ({row_reg, col_reg}<16'b0100110011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110011010001) && ({row_reg, col_reg}<16'b0100110011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110011110000) && ({row_reg, col_reg}<16'b0100110011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110011110010) && ({row_reg, col_reg}<16'b0100110011110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100110011110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110011110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100110011110110)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==16'b0100110011110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110011111000) && ({row_reg, col_reg}<16'b0100110011111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110011111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110011111011) && ({row_reg, col_reg}<16'b0100110011111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0100110011111110) && ({row_reg, col_reg}<16'b0100110100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110100000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110100000001) && ({row_reg, col_reg}<16'b0100110100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110100000101) && ({row_reg, col_reg}<16'b0100110100000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110100000111) && ({row_reg, col_reg}<16'b0100110100001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110100001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100110100001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110100001100) && ({row_reg, col_reg}<16'b0100110100001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100110100001110) && ({row_reg, col_reg}<16'b0100110100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110100010010) && ({row_reg, col_reg}<16'b0100110100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110100100110) && ({row_reg, col_reg}<16'b0100110100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110100101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100110100101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100110100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110100101101) && ({row_reg, col_reg}<16'b0100110100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110100110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100110100110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100110100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110100110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100110100111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110100111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110100111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110100111011) && ({row_reg, col_reg}<16'b0100110100111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100110100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110100111111) && ({row_reg, col_reg}<16'b0100110101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110101000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100110101000100) && ({row_reg, col_reg}<16'b0100110101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110101000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100110101000111) && ({row_reg, col_reg}<16'b0100110101001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110101001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100110101001010) && ({row_reg, col_reg}<16'b0100110101001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100110101001101) && ({row_reg, col_reg}<16'b0100110101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100110101001111) && ({row_reg, col_reg}<16'b0100110101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100110101010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100110101010101) && ({row_reg, col_reg}<16'b0100110101010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100110101010111) && ({row_reg, col_reg}<16'b0100110101011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110101011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100110101011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110101011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100110101011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110101011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100110101011110)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0100110101011111)) color_data = 12'b100010010111;
		if(({row_reg, col_reg}==16'b0100110101100000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0100110101100001)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}>=16'b0100110101100010) && ({row_reg, col_reg}<16'b0100110101100101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100110101100101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100110101100110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100110101100111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0100110101101000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0100110101101001)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==16'b0100110101101010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0100110101101011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100110101101100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0100110101101101) && ({row_reg, col_reg}<16'b0100110101101111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100110101101111)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}>=16'b0100110101110000) && ({row_reg, col_reg}<16'b0100110101110010)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0100110101110010)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0100110101110011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100110101110100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100110101110101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100110101110110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100110101110111)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0100110101111000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0100110101111001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0100110101111010)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0100110101111011)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0100110101111100)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100110101111101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0100110101111110) && ({row_reg, col_reg}<16'b0100110110000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100110110000000)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}>=16'b0100110110000001) && ({row_reg, col_reg}<16'b0100110110000011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0100110110000011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0100110110000100)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0100110110000101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0100110110000110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100110110000111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100110110001000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100110110001001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0100110110001010)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==16'b0100110110001011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=16'b0100110110001100) && ({row_reg, col_reg}<16'b0100110110001110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100110110001110)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0100110110001111)) color_data = 12'b110011001001;
		if(({row_reg, col_reg}==16'b0100110110010000)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0100110110010001)) color_data = 12'b110011001001;
		if(({row_reg, col_reg}==16'b0100110110010010)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0100110110010011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=16'b0100110110010100) && ({row_reg, col_reg}<16'b0100110110010111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100110110010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100110110011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110110011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100110110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100110110011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100110110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100110110011101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0100110110011110) && ({row_reg, col_reg}<16'b0100110110100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100110110100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100110110100001) && ({row_reg, col_reg}<16'b0100110110100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100110110100011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100110110100100) && ({row_reg, col_reg}<16'b0100110110100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100110110100111) && ({row_reg, col_reg}<16'b0100110110101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100110110101100) && ({row_reg, col_reg}<16'b0100110110110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100110110110000) && ({row_reg, col_reg}<16'b0100110110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100110110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100110110110100) && ({row_reg, col_reg}<16'b0100110110110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100110110110110) && ({row_reg, col_reg}<16'b0100110110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100110110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100110110111001) && ({row_reg, col_reg}<16'b0100110110111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100110110111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100110110111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110110111110) && ({row_reg, col_reg}<16'b0100110111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110111000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100110111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110111000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100110111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110111000100) && ({row_reg, col_reg}<16'b0100110111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100110111000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110111000111) && ({row_reg, col_reg}<16'b0100110111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100110111001011) && ({row_reg, col_reg}<16'b0100110111001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110111001111) && ({row_reg, col_reg}<16'b0100110111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110111010001) && ({row_reg, col_reg}<16'b0100110111110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110111110000) && ({row_reg, col_reg}<16'b0100110111110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110111110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110111110110) && ({row_reg, col_reg}<16'b0100110111111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100110111111011) && ({row_reg, col_reg}<16'b0100110111111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0100110111111110) && ({row_reg, col_reg}<16'b0100111000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100111000000000) && ({row_reg, col_reg}<16'b0100111000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111000000101) && ({row_reg, col_reg}<16'b0100111000001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100111000001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111000001001) && ({row_reg, col_reg}<16'b0100111000001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111000001101) && ({row_reg, col_reg}<16'b0100111000001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111000001111) && ({row_reg, col_reg}<16'b0100111000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111000010011) && ({row_reg, col_reg}<16'b0100111000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100111000100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100111000100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111000100111) && ({row_reg, col_reg}<16'b0100111000101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100111000101001) && ({row_reg, col_reg}<16'b0100111000101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111000101110) && ({row_reg, col_reg}<16'b0100111000110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111000110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111000110010) && ({row_reg, col_reg}<16'b0100111000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111000110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100111000110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111000110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100111000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111000111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111000111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111000111011) && ({row_reg, col_reg}<16'b0100111000111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100111000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111000111111) && ({row_reg, col_reg}<16'b0100111001000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111001000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100111001000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100111001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100111001000111) && ({row_reg, col_reg}<16'b0100111001001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111001001001) && ({row_reg, col_reg}<16'b0100111001001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100111001001100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100111001001101) && ({row_reg, col_reg}<16'b0100111001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100111001001111) && ({row_reg, col_reg}<16'b0100111001010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100111001010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100111001011000) && ({row_reg, col_reg}<16'b0100111001011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100111001011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100111001011011) && ({row_reg, col_reg}<16'b0100111001011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100111001011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100111001011110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100111001011111)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0100111001100000)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0100111001100001)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0100111001100010)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0100111001100011)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0100111001100100)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0100111001100101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100111001100110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100111001100111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100111001101000)) color_data = 12'b010101100100;
		if(({row_reg, col_reg}==16'b0100111001101001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100111001101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0100111001101011) && ({row_reg, col_reg}<16'b0100111001101101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100111001101101)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0100111001101110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100111001101111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100111001110000)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0100111001110001)) color_data = 12'b010101100100;
		if(({row_reg, col_reg}==16'b0100111001110010)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100111001110011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100111001110100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0100111001110101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100111001110110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100111001110111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0100111001111000) && ({row_reg, col_reg}<16'b0100111001111011)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0100111001111011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100111001111100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100111001111101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0100111001111110)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0100111001111111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100111010000000)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}>=16'b0100111010000001) && ({row_reg, col_reg}<16'b0100111010000011)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0100111010000011)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0100111010000100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100111010000101) && ({row_reg, col_reg}<16'b0100111010000111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100111010000111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100111010001000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0100111010001001)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0100111010001010)) color_data = 12'b101111001001;
		if(({row_reg, col_reg}==16'b0100111010001011)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0100111010001100)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0100111010001101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100111010001110)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0100111010001111)) color_data = 12'b110011011010;
		if(({row_reg, col_reg}==16'b0100111010010000)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0100111010010001)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0100111010010010)) color_data = 12'b100110000110;
		if(({row_reg, col_reg}==16'b0100111010010011)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0100111010010100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100111010010101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100111010010110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100111010010111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100111010011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111010011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100111010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100111010011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100111010011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100111010011101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0100111010011110) && ({row_reg, col_reg}<16'b0100111010100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100111010100000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0100111010100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100111010100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100111010100011) && ({row_reg, col_reg}<16'b0100111010100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100111010100111) && ({row_reg, col_reg}<16'b0100111010101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100111010101100) && ({row_reg, col_reg}<16'b0100111010110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100111010110000) && ({row_reg, col_reg}<16'b0100111010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100111010110011) && ({row_reg, col_reg}<16'b0100111010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100111010110110) && ({row_reg, col_reg}<16'b0100111010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100111010111000) && ({row_reg, col_reg}<16'b0100111010111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111010111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100111010111100) && ({row_reg, col_reg}<16'b0100111011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111011000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100111011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111011000100) && ({row_reg, col_reg}<16'b0100111011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111011000110) && ({row_reg, col_reg}<16'b0100111011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111011001000) && ({row_reg, col_reg}<16'b0100111011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100111011001010) && ({row_reg, col_reg}<16'b0100111011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111011010001) && ({row_reg, col_reg}<16'b0100111011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111011110000) && ({row_reg, col_reg}<16'b0100111011110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111011110100) && ({row_reg, col_reg}<16'b0100111011110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111011110110) && ({row_reg, col_reg}<16'b0100111011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100111011111001) && ({row_reg, col_reg}<16'b0100111011111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111011111011) && ({row_reg, col_reg}<16'b0100111011111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0100111011111110) && ({row_reg, col_reg}<16'b0100111100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100111100000000) && ({row_reg, col_reg}<16'b0100111100000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111100000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100111100000011) && ({row_reg, col_reg}<16'b0100111100001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111100001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111100001101) && ({row_reg, col_reg}<16'b0100111100001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100111100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111100010000) && ({row_reg, col_reg}<16'b0100111100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111100010011) && ({row_reg, col_reg}<16'b0100111100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111100100100) && ({row_reg, col_reg}<16'b0100111100100110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111100100110) && ({row_reg, col_reg}<16'b0100111100101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100111100101001) && ({row_reg, col_reg}<16'b0100111100101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111100101110) && ({row_reg, col_reg}<16'b0100111100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111100110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111100110010) && ({row_reg, col_reg}<16'b0100111100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111100110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100111100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111100110111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100111100111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100111100111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100111100111010) && ({row_reg, col_reg}<16'b0100111100111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111100111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100111100111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100111100111110) && ({row_reg, col_reg}<16'b0100111101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111101000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100111101000100) && ({row_reg, col_reg}<16'b0100111101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100111101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111101000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100111101001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111101001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100111101001010) && ({row_reg, col_reg}<16'b0100111101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100111101001100) && ({row_reg, col_reg}<16'b0100111101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100111101001111) && ({row_reg, col_reg}<16'b0100111101010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100111101010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100111101010011) && ({row_reg, col_reg}<16'b0100111101010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100111101010111) && ({row_reg, col_reg}<16'b0100111101011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100111101011010) && ({row_reg, col_reg}<16'b0100111101011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100111101011100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0100111101011101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0100111101011110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100111101011111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0100111101100000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100111101100001)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==16'b0100111101100010)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0100111101100011)) color_data = 12'b110111011011;
		if(({row_reg, col_reg}==16'b0100111101100100)) color_data = 12'b101110111000;
		if(({row_reg, col_reg}==16'b0100111101100101)) color_data = 12'b011001110101;
		if(({row_reg, col_reg}>=16'b0100111101100110) && ({row_reg, col_reg}<16'b0100111101101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100111101101000) && ({row_reg, col_reg}<16'b0100111101101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111101101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100111101101100) && ({row_reg, col_reg}<16'b0100111101101111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100111101101111)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0100111101110000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100111101110001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100111101110010)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}>=16'b0100111101110011) && ({row_reg, col_reg}<16'b0100111101110110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100111101110110) && ({row_reg, col_reg}<16'b0100111101111101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100111101111101) && ({row_reg, col_reg}<16'b0100111101111111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100111101111111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100111110000000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100111110000001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0100111110000010) && ({row_reg, col_reg}<16'b0100111110000111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100111110000111)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0100111110001000)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0100111110001001)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0100111110001010)) color_data = 12'b110010111001;
		if(({row_reg, col_reg}==16'b0100111110001011)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0100111110001100)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0100111110001101)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100111110001110)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0100111110001111)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0100111110010000)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0100111110010001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0100111110010010) && ({row_reg, col_reg}<16'b0100111110010100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100111110010100)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100111110010101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100111110010110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100111110010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100111110011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111110011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100111110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100111110011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100111110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100111110011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100111110011110) && ({row_reg, col_reg}<16'b0100111110100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100111110100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100111110100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100111110100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100111110100011) && ({row_reg, col_reg}<16'b0100111110100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100111110100111) && ({row_reg, col_reg}<16'b0100111110101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100111110101100) && ({row_reg, col_reg}<16'b0100111110110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100111110110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100111110110001) && ({row_reg, col_reg}<16'b0100111110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100111110110100) && ({row_reg, col_reg}<16'b0100111110110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100111110110110) && ({row_reg, col_reg}<16'b0100111110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100111110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100111110111001) && ({row_reg, col_reg}<16'b0100111110111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100111110111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100111110111101) && ({row_reg, col_reg}<16'b0100111110111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100111110111111) && ({row_reg, col_reg}<16'b0100111111000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111111000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100111111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111111000100) && ({row_reg, col_reg}<16'b0100111111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111111000110) && ({row_reg, col_reg}<16'b0100111111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111111001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100111111001010) && ({row_reg, col_reg}<16'b0100111111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111111010001) && ({row_reg, col_reg}<16'b0100111111110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100111111110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100111111110001) && ({row_reg, col_reg}<16'b0100111111110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111111110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100111111110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111111110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111111111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100111111111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111111111011) && ({row_reg, col_reg}<16'b0100111111111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0100111111111110) && ({row_reg, col_reg}<16'b0101000000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000000000001) && ({row_reg, col_reg}<16'b0101000000000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101000000000100) && ({row_reg, col_reg}<16'b0101000000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000000001101) && ({row_reg, col_reg}<16'b0101000000001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101000000001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000000010000) && ({row_reg, col_reg}<16'b0101000000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000000010011) && ({row_reg, col_reg}<16'b0101000000100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101000000100100) && ({row_reg, col_reg}<16'b0101000000100110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000000100110) && ({row_reg, col_reg}<16'b0101000000101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000000101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000000101001) && ({row_reg, col_reg}<16'b0101000000101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000000101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101000000101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000000101110) && ({row_reg, col_reg}<16'b0101000000110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000000110000) && ({row_reg, col_reg}<16'b0101000000110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000000110010) && ({row_reg, col_reg}<16'b0101000000110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000000110111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0101000000111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101000000111001) && ({row_reg, col_reg}<16'b0101000000111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101000000111011) && ({row_reg, col_reg}<16'b0101000001000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000001000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000001000100) && ({row_reg, col_reg}<16'b0101000001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000001000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101000001000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000001001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101000001001001) && ({row_reg, col_reg}<16'b0101000001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101000001001100) && ({row_reg, col_reg}<16'b0101000001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000001001111) && ({row_reg, col_reg}<16'b0101000001010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101000001010111) && ({row_reg, col_reg}<16'b0101000001011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000001011001) && ({row_reg, col_reg}<16'b0101000001011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000001011100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0101000001011101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0101000001011110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101000001011111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101000001100000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101000001100001)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0101000001100010)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0101000001100011)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==16'b0101000001100100)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0101000001100101)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0101000001100110)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0101000001100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000001101000) && ({row_reg, col_reg}<16'b0101000001101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000001101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000001101011) && ({row_reg, col_reg}<16'b0101000001101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000001101101) && ({row_reg, col_reg}<16'b0101000001101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000001101111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0101000001110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101000001110001) && ({row_reg, col_reg}<16'b0101000001110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101000001110011) && ({row_reg, col_reg}<16'b0101000001110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101000001110111) && ({row_reg, col_reg}<16'b0101000001111101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0101000001111101) && ({row_reg, col_reg}<16'b0101000001111111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101000001111111)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0101000010000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101000010000001) && ({row_reg, col_reg}<16'b0101000010000011)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0101000010000011) && ({row_reg, col_reg}<16'b0101000010000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101000010000101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101000010000110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101000010000111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0101000010001000)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0101000010001001)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==16'b0101000010001010)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0101000010001011)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==16'b0101000010001100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101000010001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101000010001110)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0101000010001111)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0101000010010000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101000010010001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0101000010010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101000010010011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101000010010100)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0101000010010101)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0101000010010110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101000010010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101000010011000) && ({row_reg, col_reg}<16'b0101000010011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101000010011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101000010011100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101000010011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101000010011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000010011111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0101000010100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101000010100001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101000010100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101000010100011) && ({row_reg, col_reg}<16'b0101000010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101000010100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0101000010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000010101001) && ({row_reg, col_reg}<16'b0101000010101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000010101011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101000010101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101000010101101) && ({row_reg, col_reg}<16'b0101000010110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101000010110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101000010110001) && ({row_reg, col_reg}<16'b0101000010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000010110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101000010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000010110110) && ({row_reg, col_reg}<16'b0101000010111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101000010111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000010111101) && ({row_reg, col_reg}<16'b0101000010111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101000010111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101000011000000) && ({row_reg, col_reg}<16'b0101000011000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000011000010) && ({row_reg, col_reg}<16'b0101000011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101000011000100) && ({row_reg, col_reg}<16'b0101000011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000011000110) && ({row_reg, col_reg}<16'b0101000011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000011001001) && ({row_reg, col_reg}<16'b0101000011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000011001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000011001100) && ({row_reg, col_reg}<16'b0101000011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000011010001) && ({row_reg, col_reg}<16'b0101000011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101000011110000) && ({row_reg, col_reg}<16'b0101000011110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000011110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000011110011) && ({row_reg, col_reg}<16'b0101000011111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000011111000) && ({row_reg, col_reg}<16'b0101000011111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000011111011) && ({row_reg, col_reg}<16'b0101000011111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0101000011111110) && ({row_reg, col_reg}<16'b0101000100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000100000001) && ({row_reg, col_reg}<16'b0101000100000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101000100000101) && ({row_reg, col_reg}<16'b0101000100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000100001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101000100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101000100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000100010000) && ({row_reg, col_reg}<16'b0101000100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000100010010) && ({row_reg, col_reg}<16'b0101000100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101000100100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000100100110) && ({row_reg, col_reg}<16'b0101000100101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000100101001) && ({row_reg, col_reg}<16'b0101000100101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000100101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101000100101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000100101110) && ({row_reg, col_reg}<16'b0101000100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000100110000) && ({row_reg, col_reg}<16'b0101000100110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000100110010) && ({row_reg, col_reg}<16'b0101000100110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000100110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101000100111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101000100111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101000100111010) && ({row_reg, col_reg}<16'b0101000101000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000101000010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101000101000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000101000100) && ({row_reg, col_reg}<16'b0101000101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101000101000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000101001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101000101001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000101001010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101000101001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101000101001100) && ({row_reg, col_reg}<16'b0101000101001110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0101000101001110) && ({row_reg, col_reg}<16'b0101000101010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101000101010110) && ({row_reg, col_reg}<16'b0101000101011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000101011010) && ({row_reg, col_reg}<16'b0101000101011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000101011100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0101000101011101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0101000101011110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101000101011111)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0101000101100000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101000101100001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101000101100010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=16'b0101000101100011) && ({row_reg, col_reg}<16'b0101000101100101)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0101000101100101)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0101000101100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101000101100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000101101000) && ({row_reg, col_reg}<16'b0101000101101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101000101101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101000101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000101101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000101101101) && ({row_reg, col_reg}<16'b0101000101110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000101110001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101000101110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000101110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101000101110100) && ({row_reg, col_reg}<16'b0101000101110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101000101110111)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0101000101111000) && ({row_reg, col_reg}<16'b0101000110000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101000110000101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0101000110000110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101000110000111)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=16'b0101000110001000) && ({row_reg, col_reg}<16'b0101000110001010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0101000110001010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101000110001011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101000110001100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101000110001101)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0101000110001110) && ({row_reg, col_reg}<16'b0101000110010001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101000110010001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101000110010010) && ({row_reg, col_reg}<16'b0101000110010100)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0101000110010100) && ({row_reg, col_reg}<16'b0101000110010110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101000110010110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101000110010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101000110011000) && ({row_reg, col_reg}<16'b0101000110011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101000110011011) && ({row_reg, col_reg}<16'b0101000110011101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101000110011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101000110011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101000110011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000110100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101000110100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101000110100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101000110100011) && ({row_reg, col_reg}<16'b0101000110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101000110100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0101000110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000110101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000110101010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0101000110101011) && ({row_reg, col_reg}<16'b0101000110101101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0101000110101101) && ({row_reg, col_reg}<16'b0101000110101111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101000110101111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101000110110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000110110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000110110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101000110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000110110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101000110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000110110110) && ({row_reg, col_reg}<16'b0101000110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101000110111000) && ({row_reg, col_reg}<16'b0101000110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000110111010) && ({row_reg, col_reg}<16'b0101000110111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101000110111100) && ({row_reg, col_reg}<16'b0101000110111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101000110111110) && ({row_reg, col_reg}<16'b0101000111000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101000111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000111000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101000111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101000111000100) && ({row_reg, col_reg}<16'b0101000111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000111000110) && ({row_reg, col_reg}<16'b0101000111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000111001001) && ({row_reg, col_reg}<16'b0101000111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000111001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000111001100) && ({row_reg, col_reg}<16'b0101000111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000111010001) && ({row_reg, col_reg}<16'b0101000111110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101000111110000) && ({row_reg, col_reg}<16'b0101000111110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000111110011) && ({row_reg, col_reg}<16'b0101000111110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000111110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101000111111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101000111111001) && ({row_reg, col_reg}<16'b0101000111111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000111111011) && ({row_reg, col_reg}<16'b0101000111111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101000111111110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0101000111111111) && ({row_reg, col_reg}<16'b0101001000000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001000000010) && ({row_reg, col_reg}<16'b0101001000001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101001000001000) && ({row_reg, col_reg}<16'b0101001000001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001000001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001000001111) && ({row_reg, col_reg}<16'b0101001000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001000010010) && ({row_reg, col_reg}<16'b0101001000100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101001000100110) && ({row_reg, col_reg}<16'b0101001000101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101001000101001) && ({row_reg, col_reg}<16'b0101001000101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001000101110) && ({row_reg, col_reg}<16'b0101001000110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101001000110000) && ({row_reg, col_reg}<16'b0101001000110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001000110010) && ({row_reg, col_reg}<16'b0101001000110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001000110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101001000110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101001000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001000110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001000111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101001000111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101001000111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001000111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001000111100) && ({row_reg, col_reg}<16'b0101001000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101001000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001000111111) && ({row_reg, col_reg}<16'b0101001001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001001000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101001001000010) && ({row_reg, col_reg}<16'b0101001001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001001000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101001001000111) && ({row_reg, col_reg}<16'b0101001001001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101001001001001) && ({row_reg, col_reg}<16'b0101001001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101001001001100) && ({row_reg, col_reg}<16'b0101001001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101001001001111) && ({row_reg, col_reg}<16'b0101001001010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101001001010111) && ({row_reg, col_reg}<16'b0101001001011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001001011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101001001011100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0101001001011101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0101001001011110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101001001011111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101001001100000) && ({row_reg, col_reg}<16'b0101001001100011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101001001100011)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0101001001100100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101001001100101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101001001100110)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0101001001100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101001001101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001001101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101001001101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001001101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101001001101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101001001101101) && ({row_reg, col_reg}<16'b0101001001101111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001001101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101001001110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001001110001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101001001110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001001110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101001001110100) && ({row_reg, col_reg}<16'b0101001001110110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101001001110110) && ({row_reg, col_reg}<16'b0101001001111000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101001001111000)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0101001001111001) && ({row_reg, col_reg}<16'b0101001010000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001010000101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101001010000110)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0101001010000111) && ({row_reg, col_reg}<16'b0101001010001001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101001010001001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101001010001010)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0101001010001011) && ({row_reg, col_reg}<16'b0101001010001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101001010001101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0101001010001110) && ({row_reg, col_reg}<16'b0101001010010001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101001010010001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101001010010010)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0101001010010011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101001010010100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101001010010101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101001010010110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101001010010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101001010011000) && ({row_reg, col_reg}<16'b0101001010011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101001010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101001010011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101001010011100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101001010011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001010011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001010011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101001010100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0101001010100001) && ({row_reg, col_reg}<16'b0101001010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101001010100011) && ({row_reg, col_reg}<16'b0101001010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001010100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0101001010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101001010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001010101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101001010101010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0101001010101011) && ({row_reg, col_reg}<16'b0101001010101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101001010101101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101001010101110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101001010101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101001010110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101001010110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001010110010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0101001010110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101001010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101001010110110) && ({row_reg, col_reg}<16'b0101001010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101001010111000) && ({row_reg, col_reg}<16'b0101001010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101001010111010) && ({row_reg, col_reg}<16'b0101001010111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101001010111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101001010111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101001010111110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0101001010111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001011000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101001011000001) && ({row_reg, col_reg}<16'b0101001011000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001011000011) && ({row_reg, col_reg}<16'b0101001011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001011000110) && ({row_reg, col_reg}<16'b0101001011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001011010001) && ({row_reg, col_reg}<16'b0101001011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101001011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001011110000) && ({row_reg, col_reg}<16'b0101001011110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101001011110011) && ({row_reg, col_reg}<16'b0101001011110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001011110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101001011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101001011111001) && ({row_reg, col_reg}<16'b0101001011111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001011111011) && ({row_reg, col_reg}<16'b0101001011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101001011111110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0101001011111111) && ({row_reg, col_reg}<16'b0101001100000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001100000011) && ({row_reg, col_reg}<16'b0101001100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101001100001000) && ({row_reg, col_reg}<16'b0101001100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001100001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101001100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101001100001111) && ({row_reg, col_reg}<16'b0101001100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001100010010) && ({row_reg, col_reg}<16'b0101001100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101001100100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001100100110) && ({row_reg, col_reg}<16'b0101001100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101001100101001) && ({row_reg, col_reg}<16'b0101001100101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001100101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101001100101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001100101110) && ({row_reg, col_reg}<16'b0101001100110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001100110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001100110010) && ({row_reg, col_reg}<16'b0101001100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001100110100) && ({row_reg, col_reg}<16'b0101001100110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101001100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001100110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101001100111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001100111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101001100111010) && ({row_reg, col_reg}<16'b0101001100111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001100111100) && ({row_reg, col_reg}<16'b0101001100111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101001100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001100111111) && ({row_reg, col_reg}<16'b0101001101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001101000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101001101000010) && ({row_reg, col_reg}<16'b0101001101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101001101000100) && ({row_reg, col_reg}<16'b0101001101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101001101000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101001101000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001101001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101001101001001) && ({row_reg, col_reg}<16'b0101001101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101001101001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001101001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101001101001110) && ({row_reg, col_reg}<16'b0101001101010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101001101010000) && ({row_reg, col_reg}<16'b0101001101010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101001101010110) && ({row_reg, col_reg}<16'b0101001101011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001101011001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0101001101011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001101011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101001101011100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0101001101011101) && ({row_reg, col_reg}<16'b0101001101011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101001101011111) && ({row_reg, col_reg}<16'b0101001101100001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101001101100001) && ({row_reg, col_reg}<16'b0101001101100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101001101100100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101001101100101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0101001101100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001101100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101001101101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001101101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101001101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001101101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101001101101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101001101101101) && ({row_reg, col_reg}<16'b0101001101110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001101110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001101110001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101001101110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001101110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101001101110100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001101110101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0101001101110110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101001101110111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0101001101111000) && ({row_reg, col_reg}<16'b0101001110000111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101001110000111)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101001110001000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101001110001001) && ({row_reg, col_reg}<16'b0101001110001111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101001110001111) && ({row_reg, col_reg}<16'b0101001110010001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101001110010001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101001110010010) && ({row_reg, col_reg}<16'b0101001110010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001110010100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101001110010101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101001110010110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101001110010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101001110011000) && ({row_reg, col_reg}<16'b0101001110011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101001110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101001110011011) && ({row_reg, col_reg}<16'b0101001110011101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101001110011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101001110011110) && ({row_reg, col_reg}<16'b0101001110100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101001110100000) && ({row_reg, col_reg}<16'b0101001110100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101001110100011) && ({row_reg, col_reg}<16'b0101001110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001110100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0101001110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101001110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001110101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101001110101010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0101001110101011) && ({row_reg, col_reg}<16'b0101001110101101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101001110101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101001110101110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101001110101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101001110110000) && ({row_reg, col_reg}<16'b0101001110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101001110110011) && ({row_reg, col_reg}<16'b0101001110110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001110110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101001110111000) && ({row_reg, col_reg}<16'b0101001110111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001110111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001110111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101001110111101) && ({row_reg, col_reg}<16'b0101001111000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101001111000001) && ({row_reg, col_reg}<16'b0101001111000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001111000011) && ({row_reg, col_reg}<16'b0101001111000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001111000101) && ({row_reg, col_reg}<16'b0101001111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001111001001) && ({row_reg, col_reg}<16'b0101001111001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001111001110) && ({row_reg, col_reg}<16'b0101001111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001111010001) && ({row_reg, col_reg}<16'b0101001111101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101001111101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101001111110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001111110001) && ({row_reg, col_reg}<16'b0101001111110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101001111110011) && ({row_reg, col_reg}<16'b0101001111111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001111111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101001111111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001111111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001111111100) && ({row_reg, col_reg}<16'b0101001111111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0101001111111110) && ({row_reg, col_reg}<16'b0101010000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010000000000) && ({row_reg, col_reg}<16'b0101010000001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101010000001000) && ({row_reg, col_reg}<16'b0101010000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010000001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101010000001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101010000001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101010000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010000010010) && ({row_reg, col_reg}<16'b0101010000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101010000100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010000100110) && ({row_reg, col_reg}<16'b0101010000101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010000101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010000101001) && ({row_reg, col_reg}<16'b0101010000101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010000101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101010000101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010000101110) && ({row_reg, col_reg}<16'b0101010000110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010000110001) && ({row_reg, col_reg}<16'b0101010000110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010000110011) && ({row_reg, col_reg}<16'b0101010000110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101010000110110) && ({row_reg, col_reg}<16'b0101010000111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010000111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101010000111010) && ({row_reg, col_reg}<16'b0101010000111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010000111111) && ({row_reg, col_reg}<16'b0101010001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010001000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101010001000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101010001000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101010001000100) && ({row_reg, col_reg}<16'b0101010001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101010001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101010001000111) && ({row_reg, col_reg}<16'b0101010001001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101010001001001) && ({row_reg, col_reg}<16'b0101010001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101010001001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101010001001101) && ({row_reg, col_reg}<16'b0101010001001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101010001010000) && ({row_reg, col_reg}<16'b0101010001010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101010001010111) && ({row_reg, col_reg}<16'b0101010001011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101010001011010) && ({row_reg, col_reg}<16'b0101010001011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101010001011101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0101010001011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101010001011111) && ({row_reg, col_reg}<16'b0101010001100001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101010001100001) && ({row_reg, col_reg}<16'b0101010001100011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101010001100011)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}>=16'b0101010001100100) && ({row_reg, col_reg}<16'b0101010001100110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101010001100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101010001100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101010001101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010001101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010001101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010001101011) && ({row_reg, col_reg}<16'b0101010001101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101010001101101) && ({row_reg, col_reg}<16'b0101010001110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101010001110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010001110001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101010001110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010001110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101010001110100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101010001110101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0101010001110110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101010001110111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101010001111000) && ({row_reg, col_reg}<16'b0101010010000110)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0101010010000110) && ({row_reg, col_reg}<16'b0101010010001010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101010010001010) && ({row_reg, col_reg}<16'b0101010010001100)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0101010010001100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101010010001101) && ({row_reg, col_reg}<16'b0101010010010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101010010010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010010010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101010010010101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101010010010110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101010010010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101010010011000) && ({row_reg, col_reg}<16'b0101010010011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101010010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101010010011011) && ({row_reg, col_reg}<16'b0101010010011101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101010010011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101010010011110) && ({row_reg, col_reg}<16'b0101010010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101010010100011) && ({row_reg, col_reg}<16'b0101010010100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101010010100111) && ({row_reg, col_reg}<16'b0101010010110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101010010110001) && ({row_reg, col_reg}<16'b0101010010110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101010010110111) && ({row_reg, col_reg}<16'b0101010010111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101010010111010) && ({row_reg, col_reg}<16'b0101010010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010010111101) && ({row_reg, col_reg}<16'b0101010011000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101010011000001) && ({row_reg, col_reg}<16'b0101010011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010011001001) && ({row_reg, col_reg}<16'b0101010011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101010011001011) && ({row_reg, col_reg}<16'b0101010011001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010011001111) && ({row_reg, col_reg}<16'b0101010011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010011010001) && ({row_reg, col_reg}<16'b0101010011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101010011110000) && ({row_reg, col_reg}<16'b0101010011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101010011110011) && ({row_reg, col_reg}<16'b0101010011110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010011110101) && ({row_reg, col_reg}<16'b0101010011110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010011110111) && ({row_reg, col_reg}<16'b0101010011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010011111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101010011111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010011111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010011111100) && ({row_reg, col_reg}<16'b0101010011111110)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0101010011111110) && ({row_reg, col_reg}<16'b0101010100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010100000000) && ({row_reg, col_reg}<16'b0101010100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101010100001000) && ({row_reg, col_reg}<16'b0101010100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010100001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101010100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101010100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101010100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010100010010) && ({row_reg, col_reg}<16'b0101010100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101010100100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010100100110) && ({row_reg, col_reg}<16'b0101010100101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010100101001) && ({row_reg, col_reg}<16'b0101010100101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010100101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101010100101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010100101110) && ({row_reg, col_reg}<16'b0101010100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010100110000) && ({row_reg, col_reg}<16'b0101010100110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010100110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101010100110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101010100110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010100110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101010100111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010100111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101010100111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010100111011) && ({row_reg, col_reg}<16'b0101010101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010101000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101010101000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101010101000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010101000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101010101000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101010101000110) && ({row_reg, col_reg}<16'b0101010101001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101010101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101010101001010) && ({row_reg, col_reg}<16'b0101010101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101010101001100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101010101001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010101001110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101010101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101010101010000) && ({row_reg, col_reg}<16'b0101010101011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101010101011000) && ({row_reg, col_reg}<16'b0101010101011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101010101011010) && ({row_reg, col_reg}<16'b0101010101011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101010101011101) && ({row_reg, col_reg}<16'b0101010101100000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101010101100000) && ({row_reg, col_reg}<16'b0101010101100011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101010101100011)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0101010101100100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101010101100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101010101100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101010101100111) && ({row_reg, col_reg}<16'b0101010101101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101010101101101) && ({row_reg, col_reg}<16'b0101010101110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101010101110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010101110001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101010101110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010101110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101010101110100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101010101110101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0101010101110110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101010101110111) && ({row_reg, col_reg}<16'b0101010110000111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101010110000111)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0101010110001000)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0101010110001001) && ({row_reg, col_reg}<16'b0101010110001011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101010110001011)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0101010110001100) && ({row_reg, col_reg}<16'b0101010110010011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101010110010011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==16'b0101010110010100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101010110010101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101010110010110)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0101010110010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101010110011000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101010110011001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101010110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101010110011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101010110011100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101010110011101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0101010110011110) && ({row_reg, col_reg}<16'b0101010110100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101010110100011) && ({row_reg, col_reg}<16'b0101010110100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101010110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101010110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101010110101001) && ({row_reg, col_reg}<16'b0101010110110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101010110110000) && ({row_reg, col_reg}<16'b0101010110110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010110110010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0101010110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101010110110100) && ({row_reg, col_reg}<16'b0101010110110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010110110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101010110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010110111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101010110111010) && ({row_reg, col_reg}<16'b0101010110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010110111101) && ({row_reg, col_reg}<16'b0101010110111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101010110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101010111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010111000001) && ({row_reg, col_reg}<16'b0101010111000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010111000011) && ({row_reg, col_reg}<16'b0101010111000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010111000101) && ({row_reg, col_reg}<16'b0101010111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010111001000) && ({row_reg, col_reg}<16'b0101010111001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010111001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101010111001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010111001100) && ({row_reg, col_reg}<16'b0101010111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010111001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010111001111) && ({row_reg, col_reg}<16'b0101010111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010111010001) && ({row_reg, col_reg}<16'b0101010111101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101010111101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101010111110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010111110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101010111110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101010111110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010111110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101010111110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010111110111) && ({row_reg, col_reg}<16'b0101010111111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010111111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010111111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101010111111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010111111110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0101010111111111) && ({row_reg, col_reg}<16'b0101011000000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011000000001) && ({row_reg, col_reg}<16'b0101011000001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101011000001000) && ({row_reg, col_reg}<16'b0101011000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011000001101) && ({row_reg, col_reg}<16'b0101011000010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101011000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011000010010) && ({row_reg, col_reg}<16'b0101011000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101011000100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101011000100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011000100111) && ({row_reg, col_reg}<16'b0101011000101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011000101001) && ({row_reg, col_reg}<16'b0101011000101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011000101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101011000101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011000101110) && ({row_reg, col_reg}<16'b0101011000110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011000110000) && ({row_reg, col_reg}<16'b0101011000110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011000110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101011000110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101011000110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101011000110101) && ({row_reg, col_reg}<16'b0101011000110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101011000110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101011000111000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0101011000111001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0101011000111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011000111011) && ({row_reg, col_reg}<16'b0101011001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101011001000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101011001000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101011001000011) && ({row_reg, col_reg}<16'b0101011001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011001000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101011001000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011001001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101011001001001) && ({row_reg, col_reg}<16'b0101011001001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101011001001100) && ({row_reg, col_reg}<16'b0101011001001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101011001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101011001001111) && ({row_reg, col_reg}<16'b0101011001011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101011001011101) && ({row_reg, col_reg}<16'b0101011001011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101011001011111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101011001100000)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0101011001100001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101011001100010)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0101011001100011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101011001100100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101011001100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101011001100110) && ({row_reg, col_reg}<16'b0101011001101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011001101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101011001101001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101011001101010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0101011001101011) && ({row_reg, col_reg}<16'b0101011001101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101011001101101) && ({row_reg, col_reg}<16'b0101011001110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101011001110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011001110001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101011001110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011001110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101011001110100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101011001110101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0101011001110110) && ({row_reg, col_reg}<16'b0101011010001100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101011010001100) && ({row_reg, col_reg}<16'b0101011010001110)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0101011010001110) && ({row_reg, col_reg}<16'b0101011010010000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101011010010000)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0101011010010001) && ({row_reg, col_reg}<16'b0101011010010011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101011010010011)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0101011010010100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101011010010101)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0101011010010110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011010010111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101011010011000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101011010011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101011010011010) && ({row_reg, col_reg}<16'b0101011010011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101011010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101011010011101) && ({row_reg, col_reg}<16'b0101011010100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101011010100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0101011010100001) && ({row_reg, col_reg}<16'b0101011010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101011010100011) && ({row_reg, col_reg}<16'b0101011010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101011010100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0101011010100111) && ({row_reg, col_reg}<16'b0101011010110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101011010110000) && ({row_reg, col_reg}<16'b0101011010110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101011010110010) && ({row_reg, col_reg}<16'b0101011010110100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101011010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101011010110110) && ({row_reg, col_reg}<16'b0101011010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101011010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011010111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101011010111010)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b0101011010111011) && ({row_reg, col_reg}<16'b0101011010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101011010111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101011010111110) && ({row_reg, col_reg}<16'b0101011011000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011011000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101011011000001) && ({row_reg, col_reg}<16'b0101011011000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011011000100) && ({row_reg, col_reg}<16'b0101011011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101011011001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011011001100) && ({row_reg, col_reg}<16'b0101011011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011011001111) && ({row_reg, col_reg}<16'b0101011011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011011010001) && ({row_reg, col_reg}<16'b0101011011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101011011101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101011011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011011110001) && ({row_reg, col_reg}<16'b0101011011110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101011011110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101011011110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011011110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011011110110) && ({row_reg, col_reg}<16'b0101011011111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011011111010) && ({row_reg, col_reg}<16'b0101011011111110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0101011011111110) && ({row_reg, col_reg}<16'b0101011100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011100000000) && ({row_reg, col_reg}<16'b0101011100000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011100000010) && ({row_reg, col_reg}<16'b0101011100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101011100001000) && ({row_reg, col_reg}<16'b0101011100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011100001101) && ({row_reg, col_reg}<16'b0101011100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011100001111) && ({row_reg, col_reg}<16'b0101011100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011100010010) && ({row_reg, col_reg}<16'b0101011100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101011100100100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101011100100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011100100110) && ({row_reg, col_reg}<16'b0101011100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011100101000) && ({row_reg, col_reg}<16'b0101011100101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011100101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101011100101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011100101110) && ({row_reg, col_reg}<16'b0101011100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101011100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011100110001) && ({row_reg, col_reg}<16'b0101011100110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101011100110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011100110100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101011100110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101011100110110) && ({row_reg, col_reg}<16'b0101011100111000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101011100111000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0101011100111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101011100111010) && ({row_reg, col_reg}<16'b0101011100111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011100111100) && ({row_reg, col_reg}<16'b0101011101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101011101000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101011101000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101011101000011) && ({row_reg, col_reg}<16'b0101011101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101011101000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011101001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101011101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101011101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011101001100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101011101001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101011101001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011101001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101011101010000) && ({row_reg, col_reg}<16'b0101011101010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0101011101010011) && ({row_reg, col_reg}<16'b0101011101011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101011101011100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0101011101011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101011101011110) && ({row_reg, col_reg}<16'b0101011101100001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101011101100001) && ({row_reg, col_reg}<16'b0101011101100011)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0101011101100011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101011101100100) && ({row_reg, col_reg}<16'b0101011101100110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101011101100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101011101100111) && ({row_reg, col_reg}<16'b0101011101101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101011101101001) && ({row_reg, col_reg}<16'b0101011101101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101011101101011) && ({row_reg, col_reg}<16'b0101011101101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101011101101101) && ({row_reg, col_reg}<16'b0101011101110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101011101110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101011101110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101011101110010) && ({row_reg, col_reg}<16'b0101011101110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101011101110100) && ({row_reg, col_reg}<16'b0101011101110110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101011101110110) && ({row_reg, col_reg}<16'b0101011110001000)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0101011110001000) && ({row_reg, col_reg}<16'b0101011110001010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101011110001010)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0101011110001011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101011110001100)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0101011110001101) && ({row_reg, col_reg}<16'b0101011110001111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101011110001111)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0101011110010000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101011110010001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101011110010010)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0101011110010011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101011110010100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101011110010101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0101011110010110)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0101011110010111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101011110011000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101011110011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101011110011010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101011110011011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011110011100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0101011110011101) && ({row_reg, col_reg}<16'b0101011110100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101011110100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0101011110100001) && ({row_reg, col_reg}<16'b0101011110100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101011110100011) && ({row_reg, col_reg}<16'b0101011110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101011110100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0101011110100111) && ({row_reg, col_reg}<16'b0101011110101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101011110101011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101011110101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101011110101101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0101011110101110) && ({row_reg, col_reg}<16'b0101011110110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101011110110000) && ({row_reg, col_reg}<16'b0101011110110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011110110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101011110110011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0101011110110100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0101011110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101011110110110) && ({row_reg, col_reg}<16'b0101011110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101011110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101011110111001) && ({row_reg, col_reg}<16'b0101011110111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101011110111100) && ({row_reg, col_reg}<16'b0101011110111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101011110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011110111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101011111000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101011111000001) && ({row_reg, col_reg}<16'b0101011111000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101011111000011) && ({row_reg, col_reg}<16'b0101011111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101011111001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011111001100) && ({row_reg, col_reg}<16'b0101011111001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011111001111) && ({row_reg, col_reg}<16'b0101011111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011111010001) && ({row_reg, col_reg}<16'b0101011111101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101011111101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101011111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011111110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101011111110001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==16'b0101011111110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101011111110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101011111110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011111110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011111110110) && ({row_reg, col_reg}<16'b0101011111111001)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0101011111111001) && ({row_reg, col_reg}<16'b0101100000000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100000000001) && ({row_reg, col_reg}<16'b0101100000000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101100000000110) && ({row_reg, col_reg}<16'b0101100000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100000001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101100000001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101100000001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101100000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100000010010) && ({row_reg, col_reg}<16'b0101100000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101100000100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100000100110) && ({row_reg, col_reg}<16'b0101100000101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100000101000) && ({row_reg, col_reg}<16'b0101100000101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100000101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101100000101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100000101110) && ({row_reg, col_reg}<16'b0101100000110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100000110000) && ({row_reg, col_reg}<16'b0101100000110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100000110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101100000110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100000110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101100000110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101100000110110) && ({row_reg, col_reg}<16'b0101100000111001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101100000111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101100000111010) && ({row_reg, col_reg}<16'b0101100000111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100000111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100000111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101100000111110) && ({row_reg, col_reg}<16'b0101100001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100001000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101100001000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101100001000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101100001000100) && ({row_reg, col_reg}<16'b0101100001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101100001000110) && ({row_reg, col_reg}<16'b0101100001001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101100001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101100001001010) && ({row_reg, col_reg}<16'b0101100001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101100001001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101100001001101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101100001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100001001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101100001010000) && ({row_reg, col_reg}<16'b0101100001010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0101100001010011) && ({row_reg, col_reg}<16'b0101100001011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101100001011100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0101100001011101) && ({row_reg, col_reg}<16'b0101100001011111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101100001011111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101100001100000)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0101100001100001) && ({row_reg, col_reg}<16'b0101100001100110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101100001100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101100001100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101100001101000) && ({row_reg, col_reg}<16'b0101100001101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101100001101011) && ({row_reg, col_reg}<16'b0101100001101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101100001101101) && ({row_reg, col_reg}<16'b0101100001110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101100001110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101100001110001) && ({row_reg, col_reg}<16'b0101100001110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100001110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101100001110100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101100001110101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0101100001110110) && ({row_reg, col_reg}<16'b0101100010001001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101100010001001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101100010001010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101100010001011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101100010001100)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0101100010001101) && ({row_reg, col_reg}<16'b0101100010010001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101100010010001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0101100010010010) && ({row_reg, col_reg}<16'b0101100010010100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101100010010100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101100010010101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0101100010010110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0101100010010111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101100010011000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101100010011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101100010011010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101100010011011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101100010011100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0101100010011101) && ({row_reg, col_reg}<16'b0101100010100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101100010100000) && ({row_reg, col_reg}<16'b0101100010100010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101100010100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101100010100011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0101100010100100) && ({row_reg, col_reg}<16'b0101100010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101100010100110) && ({row_reg, col_reg}<16'b0101100010101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101100010101001) && ({row_reg, col_reg}<16'b0101100010101111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101100010101111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0101100010110000) && ({row_reg, col_reg}<16'b0101100010110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101100010110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101100010110011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0101100010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101100010110110) && ({row_reg, col_reg}<16'b0101100010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101100010111000) && ({row_reg, col_reg}<16'b0101100010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101100010111010) && ({row_reg, col_reg}<16'b0101100010111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101100010111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100010111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101100010111110) && ({row_reg, col_reg}<16'b0101100011000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100011000000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0101100011000001) && ({row_reg, col_reg}<16'b0101100011000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101100011000011) && ({row_reg, col_reg}<16'b0101100011000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100011000111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101100011001000) && ({row_reg, col_reg}<16'b0101100011001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100011001011) && ({row_reg, col_reg}<16'b0101100011001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100011001111) && ({row_reg, col_reg}<16'b0101100011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100011010001) && ({row_reg, col_reg}<16'b0101100011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101100011101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101100011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101100011110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101100011110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100011110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101100011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101100011110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100011111000) && ({row_reg, col_reg}<16'b0101100011111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100011111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100011111101) && ({row_reg, col_reg}<16'b0101100011111111)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0101100011111111) && ({row_reg, col_reg}<16'b0101100100000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101100100000110) && ({row_reg, col_reg}<16'b0101100100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100100001101) && ({row_reg, col_reg}<16'b0101100100001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101100100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101100100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100100010010) && ({row_reg, col_reg}<16'b0101100100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100100100110) && ({row_reg, col_reg}<16'b0101100100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100100101000) && ({row_reg, col_reg}<16'b0101100100101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100100101110) && ({row_reg, col_reg}<16'b0101100100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100100110000) && ({row_reg, col_reg}<16'b0101100100110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100100110010) && ({row_reg, col_reg}<16'b0101100100110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100100110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101100100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100100110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101100100111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100100111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101100100111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100100111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100100111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101100100111110) && ({row_reg, col_reg}<16'b0101100101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100101000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101100101000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101100101000011) && ({row_reg, col_reg}<16'b0101100101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100101000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101100101000111) && ({row_reg, col_reg}<16'b0101100101001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101100101001001) && ({row_reg, col_reg}<16'b0101100101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101100101001100) && ({row_reg, col_reg}<16'b0101100101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101100101001111) && ({row_reg, col_reg}<16'b0101100101010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101100101010001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0101100101010010) && ({row_reg, col_reg}<16'b0101100101010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101100101010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101100101011000) && ({row_reg, col_reg}<16'b0101100101011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101100101011100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0101100101011101) && ({row_reg, col_reg}<16'b0101100101011111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101100101011111)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0101100101100000)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0101100101100001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101100101100010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101100101100011) && ({row_reg, col_reg}<16'b0101100101100110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101100101100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101100101100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101100101101000) && ({row_reg, col_reg}<16'b0101100101101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100101101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101100101101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101100101101101) && ({row_reg, col_reg}<16'b0101100101110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101100101110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101100101110001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101100101110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100101110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101100101110100) && ({row_reg, col_reg}<16'b0101100110001001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101100110001001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101100110001010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101100110001011) && ({row_reg, col_reg}<16'b0101100110010100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101100110010100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101100110010101)) color_data = 12'b011110000110;
		if(({row_reg, col_reg}==16'b0101100110010110)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0101100110010111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101100110011000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101100110011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101100110011010) && ({row_reg, col_reg}<16'b0101100110011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101100110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101100110011101) && ({row_reg, col_reg}<16'b0101100110100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101100110100000) && ({row_reg, col_reg}<16'b0101100110100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101100110100010) && ({row_reg, col_reg}<16'b0101100110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101100110100110) && ({row_reg, col_reg}<16'b0101100110101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101100110101010) && ({row_reg, col_reg}<16'b0101100110101101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101100110101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101100110101110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101100110101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101100110110000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101100110110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101100110110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101100110110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101100110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101100110110110) && ({row_reg, col_reg}<16'b0101100110111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101100110111001) && ({row_reg, col_reg}<16'b0101100110111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100110111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101100110111100) && ({row_reg, col_reg}<16'b0101100110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101100110111111) && ({row_reg, col_reg}<16'b0101100111000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101100111000001) && ({row_reg, col_reg}<16'b0101100111000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100111000011) && ({row_reg, col_reg}<16'b0101100111000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100111000101) && ({row_reg, col_reg}<16'b0101100111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100111000111) && ({row_reg, col_reg}<16'b0101100111001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101100111001001) && ({row_reg, col_reg}<16'b0101100111001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100111001101) && ({row_reg, col_reg}<16'b0101100111001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100111001111) && ({row_reg, col_reg}<16'b0101100111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100111010001) && ({row_reg, col_reg}<16'b0101100111101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101100111101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101100111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100111110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100111110010) && ({row_reg, col_reg}<16'b0101100111110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101100111110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100111110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100111110110) && ({row_reg, col_reg}<16'b0101100111111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100111111000) && ({row_reg, col_reg}<16'b0101100111111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100111111100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0101100111111101) && ({row_reg, col_reg}<16'b0101101000000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101000000010) && ({row_reg, col_reg}<16'b0101101000000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101101000000110) && ({row_reg, col_reg}<16'b0101101000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101000001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101101000001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101101000001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101000010000) && ({row_reg, col_reg}<16'b0101101000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101000010010) && ({row_reg, col_reg}<16'b0101101000100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101101000100110) && ({row_reg, col_reg}<16'b0101101000101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101000101001) && ({row_reg, col_reg}<16'b0101101000101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101000101110) && ({row_reg, col_reg}<16'b0101101000110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101000110001) && ({row_reg, col_reg}<16'b0101101000110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101101000110011) && ({row_reg, col_reg}<16'b0101101000110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101101000110111) && ({row_reg, col_reg}<16'b0101101000111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101101000111001) && ({row_reg, col_reg}<16'b0101101000111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101000111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101101000111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101101000111110) && ({row_reg, col_reg}<16'b0101101001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101001000001) && ({row_reg, col_reg}<16'b0101101001000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101101001000100) && ({row_reg, col_reg}<16'b0101101001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101101001000110) && ({row_reg, col_reg}<16'b0101101001001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101101001001001) && ({row_reg, col_reg}<16'b0101101001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101101001001100) && ({row_reg, col_reg}<16'b0101101001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101101001001111) && ({row_reg, col_reg}<16'b0101101001010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101101001010110) && ({row_reg, col_reg}<16'b0101101001011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101101001011000) && ({row_reg, col_reg}<16'b0101101001011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101001011100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101101001011101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101101001011110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101101001011111)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0101101001100000)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0101101001100001) && ({row_reg, col_reg}<16'b0101101001100110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101101001100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101101001100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101001101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101001101001) && ({row_reg, col_reg}<16'b0101101001101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101101001101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101101001101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101101001101101) && ({row_reg, col_reg}<16'b0101101001110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101101001110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101101001110001) && ({row_reg, col_reg}<16'b0101101001110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101001110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101101001110100) && ({row_reg, col_reg}<16'b0101101001110110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101101001110110)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0101101001110111) && ({row_reg, col_reg}<16'b0101101001111100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101101001111100) && ({row_reg, col_reg}<16'b0101101001111110)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0101101001111110)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0101101001111111)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0101101010000000) && ({row_reg, col_reg}<16'b0101101010000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101101010000011) && ({row_reg, col_reg}<16'b0101101010000101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0101101010000101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0101101010000110)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0101101010000111) && ({row_reg, col_reg}<16'b0101101010001001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101101010001001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101101010001010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101101010001011) && ({row_reg, col_reg}<16'b0101101010001110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101101010001110) && ({row_reg, col_reg}<16'b0101101010010000)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0101101010010000) && ({row_reg, col_reg}<16'b0101101010010100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101101010010100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101101010010101)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0101101010010110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0101101010010111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101101010011000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101101010011001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101101010011010) && ({row_reg, col_reg}<16'b0101101010011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101101010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101101010011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101010011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101010011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101101010100000) && ({row_reg, col_reg}<16'b0101101010100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101101010100011) && ({row_reg, col_reg}<16'b0101101010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101101010100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0101101010100111) && ({row_reg, col_reg}<16'b0101101010101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101010101111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0101101010110000) && ({row_reg, col_reg}<16'b0101101010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101101010110100) && ({row_reg, col_reg}<16'b0101101010110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101101010110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101101010110111)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==16'b0101101010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101101010111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101101010111010) && ({row_reg, col_reg}<16'b0101101010111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101101010111100) && ({row_reg, col_reg}<16'b0101101010111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101010111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101101010111111) && ({row_reg, col_reg}<16'b0101101011000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101011000010) && ({row_reg, col_reg}<16'b0101101011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101011000110) && ({row_reg, col_reg}<16'b0101101011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101011001111) && ({row_reg, col_reg}<16'b0101101011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101011010001) && ({row_reg, col_reg}<16'b0101101011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101101011101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101011101111) && ({row_reg, col_reg}<16'b0101101011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101011110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101011110010) && ({row_reg, col_reg}<16'b0101101011110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101011110101) && ({row_reg, col_reg}<16'b0101101011110111)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0101101011110111) && ({row_reg, col_reg}<16'b0101101100000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101100000010) && ({row_reg, col_reg}<16'b0101101100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101101100001000) && ({row_reg, col_reg}<16'b0101101100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101100001101) && ({row_reg, col_reg}<16'b0101101100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101101100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101100010011) && ({row_reg, col_reg}<16'b0101101100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101101100100110) && ({row_reg, col_reg}<16'b0101101100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101100101001) && ({row_reg, col_reg}<16'b0101101100101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101100101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101100110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101101100110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101100110011) && ({row_reg, col_reg}<16'b0101101100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101100110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101101100110111) && ({row_reg, col_reg}<16'b0101101100111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101101100111001) && ({row_reg, col_reg}<16'b0101101100111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101100111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101101100111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101101100111110) && ({row_reg, col_reg}<16'b0101101101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101101000001) && ({row_reg, col_reg}<16'b0101101101000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101101101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101101101000111) && ({row_reg, col_reg}<16'b0101101101001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101101101001001) && ({row_reg, col_reg}<16'b0101101101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101101101001100) && ({row_reg, col_reg}<16'b0101101101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101101101001111) && ({row_reg, col_reg}<16'b0101101101010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101101101010111) && ({row_reg, col_reg}<16'b0101101101011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101101101011010) && ({row_reg, col_reg}<16'b0101101101011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101101011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101101101011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101101101011110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101101101011111)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0101101101100000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101101101100001) && ({row_reg, col_reg}<16'b0101101101100011)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0101101101100011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101101101100100) && ({row_reg, col_reg}<16'b0101101101100110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101101101100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101101101100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101101101101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101101101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101101101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101101101101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101101101101101) && ({row_reg, col_reg}<16'b0101101101110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101101101110000) && ({row_reg, col_reg}<16'b0101101101110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101101101110100) && ({row_reg, col_reg}<16'b0101101101111001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101101101111001) && ({row_reg, col_reg}<16'b0101101101111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101101101111011) && ({row_reg, col_reg}<16'b0101101110000001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101101110000001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0101101110000010) && ({row_reg, col_reg}<16'b0101101110001001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101101110001001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101101110001010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101101110001011)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0101101110001100) && ({row_reg, col_reg}<16'b0101101110001110)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101101110001110)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0101101110001111) && ({row_reg, col_reg}<16'b0101101110010100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101101110010100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101101110010101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0101101110010110)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0101101110010111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101101110011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101101110011001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0101101110011010) && ({row_reg, col_reg}<16'b0101101110011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101101110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101101110011101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0101101110011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101110011111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0101101110100000) && ({row_reg, col_reg}<16'b0101101110100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101101110100011) && ({row_reg, col_reg}<16'b0101101110100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101101110100111) && ({row_reg, col_reg}<16'b0101101110101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101110101111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0101101110110000) && ({row_reg, col_reg}<16'b0101101110110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101101110110110) && ({row_reg, col_reg}<16'b0101101110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101101110111000) && ({row_reg, col_reg}<16'b0101101110111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101101110111100) && ({row_reg, col_reg}<16'b0101101111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101111000000) && ({row_reg, col_reg}<16'b0101101111000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101111000011) && ({row_reg, col_reg}<16'b0101101111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101101111000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101111000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101111001000) && ({row_reg, col_reg}<16'b0101101111001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101111001100) && ({row_reg, col_reg}<16'b0101101111001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101111001110) && ({row_reg, col_reg}<16'b0101101111010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101111010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101111010001) && ({row_reg, col_reg}<16'b0101101111101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101101111101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101111101111) && ({row_reg, col_reg}<16'b0101101111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101111110001) && ({row_reg, col_reg}<16'b0101101111110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101111110011) && ({row_reg, col_reg}<16'b0101101111110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101111110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101111111000) && ({row_reg, col_reg}<16'b0101101111111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101111111100) && ({row_reg, col_reg}<16'b0101101111111111)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0101101111111111) && ({row_reg, col_reg}<16'b0101110000000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110000000001) && ({row_reg, col_reg}<16'b0101110000001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101110000001000) && ({row_reg, col_reg}<16'b0101110000001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110000001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101110000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110000010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101110000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110000010011) && ({row_reg, col_reg}<16'b0101110000100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101110000100110) && ({row_reg, col_reg}<16'b0101110000101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110000101010) && ({row_reg, col_reg}<16'b0101110000101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110000101110) && ({row_reg, col_reg}<16'b0101110000110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110000110000) && ({row_reg, col_reg}<16'b0101110000110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110000110010) && ({row_reg, col_reg}<16'b0101110000110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101110000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110000110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101110000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110000111001) && ({row_reg, col_reg}<16'b0101110000111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101110000111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110000111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101110000111101) && ({row_reg, col_reg}<16'b0101110001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110001000001) && ({row_reg, col_reg}<16'b0101110001000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101110001000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110001000100) && ({row_reg, col_reg}<16'b0101110001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101110001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110001000111) && ({row_reg, col_reg}<16'b0101110001001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101110001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110001001010) && ({row_reg, col_reg}<16'b0101110001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101110001001100) && ({row_reg, col_reg}<16'b0101110001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110001001111) && ({row_reg, col_reg}<16'b0101110001010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101110001010111) && ({row_reg, col_reg}<16'b0101110001011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110001011010) && ({row_reg, col_reg}<16'b0101110001011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101110001011100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101110001011101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101110001011110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101110001011111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0101110001100000) && ({row_reg, col_reg}<16'b0101110001100010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101110001100010)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0101110001100011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101110001100100) && ({row_reg, col_reg}<16'b0101110001100110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101110001100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101110001100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110001101000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==16'b0101110001101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101110001101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110001101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101110001101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110001101101) && ({row_reg, col_reg}<16'b0101110001110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101110001110000) && ({row_reg, col_reg}<16'b0101110001110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101110001110011) && ({row_reg, col_reg}<16'b0101110001110101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0101110001110101) && ({row_reg, col_reg}<16'b0101110001111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101110001111000) && ({row_reg, col_reg}<16'b0101110001111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110001111011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0101110001111100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101110001111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101110001111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110001111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101110010000000) && ({row_reg, col_reg}<16'b0101110010000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110010000010) && ({row_reg, col_reg}<16'b0101110010000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101110010000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110010000101) && ({row_reg, col_reg}<16'b0101110010000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101110010000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110010001000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101110010001001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101110010001010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101110010001011)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0101110010001100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101110010001101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101110010001110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101110010001111) && ({row_reg, col_reg}<16'b0101110010010100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101110010010100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101110010010101)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0101110010010110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101110010010111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101110010011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101110010011001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101110010011010) && ({row_reg, col_reg}<16'b0101110010011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101110010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101110010011101) && ({row_reg, col_reg}<16'b0101110010011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101110010011111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0101110010100000) && ({row_reg, col_reg}<16'b0101110010100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101110010100010) && ({row_reg, col_reg}<16'b0101110010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101110010100110) && ({row_reg, col_reg}<16'b0101110010101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101110010101011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0101110010101100) && ({row_reg, col_reg}<16'b0101110010110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101110010110000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101110010110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101110010110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101110010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101110010110100) && ({row_reg, col_reg}<16'b0101110010110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110010110110) && ({row_reg, col_reg}<16'b0101110010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101110010111000) && ({row_reg, col_reg}<16'b0101110010111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110010111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101110010111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110010111111) && ({row_reg, col_reg}<16'b0101110011000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110011000011) && ({row_reg, col_reg}<16'b0101110011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110011000110) && ({row_reg, col_reg}<16'b0101110011001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110011001100) && ({row_reg, col_reg}<16'b0101110011001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110011001110) && ({row_reg, col_reg}<16'b0101110011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110011010001) && ({row_reg, col_reg}<16'b0101110011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101110011101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101110011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110011110001) && ({row_reg, col_reg}<16'b0101110011110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110011110111) && ({row_reg, col_reg}<16'b0101110011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110011111001) && ({row_reg, col_reg}<16'b0101110011111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110011111100) && ({row_reg, col_reg}<16'b0101110011111110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0101110011111110) && ({row_reg, col_reg}<16'b0101110100000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110100000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101110100000010) && ({row_reg, col_reg}<16'b0101110100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110100000110) && ({row_reg, col_reg}<16'b0101110100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101110100001000) && ({row_reg, col_reg}<16'b0101110100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101110100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110100010011) && ({row_reg, col_reg}<16'b0101110100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101110100100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101110100100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110100100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101110100101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110100101001) && ({row_reg, col_reg}<16'b0101110100101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101110100101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110100101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101110100101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110100101110) && ({row_reg, col_reg}<16'b0101110100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110100110000) && ({row_reg, col_reg}<16'b0101110100110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110100110011) && ({row_reg, col_reg}<16'b0101110100110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101110100110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101110100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110100110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101110100111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101110100111001) && ({row_reg, col_reg}<16'b0101110100111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101110100111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110100111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101110100111110) && ({row_reg, col_reg}<16'b0101110101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110101000001) && ({row_reg, col_reg}<16'b0101110101000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101110101000011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0101110101000100) && ({row_reg, col_reg}<16'b0101110101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110101000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101110101000111) && ({row_reg, col_reg}<16'b0101110101001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101110101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110101001010) && ({row_reg, col_reg}<16'b0101110101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101110101001100) && ({row_reg, col_reg}<16'b0101110101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110101001111) && ({row_reg, col_reg}<16'b0101110101010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101110101010111) && ({row_reg, col_reg}<16'b0101110101011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110101011010) && ({row_reg, col_reg}<16'b0101110101011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101110101011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101110101011101) && ({row_reg, col_reg}<16'b0101110101011111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101110101011111)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}>=16'b0101110101100000) && ({row_reg, col_reg}<16'b0101110101100010)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0101110101100010) && ({row_reg, col_reg}<16'b0101110101100110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101110101100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101110101100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110101101000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==16'b0101110101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101110101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110101101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101110101101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110101101101) && ({row_reg, col_reg}<16'b0101110101110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101110101110000) && ({row_reg, col_reg}<16'b0101110101110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101110101110011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0101110101110100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101110101110101) && ({row_reg, col_reg}<16'b0101110101111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101110101111001) && ({row_reg, col_reg}<16'b0101110101111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110101111011) && ({row_reg, col_reg}<16'b0101110101111101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101110101111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101110101111110) && ({row_reg, col_reg}<16'b0101110110000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110110000001) && ({row_reg, col_reg}<16'b0101110110000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101110110000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101110110000101) && ({row_reg, col_reg}<16'b0101110110000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110110000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101110110001000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101110110001001) && ({row_reg, col_reg}<16'b0101110110001100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101110110001100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101110110001101) && ({row_reg, col_reg}<16'b0101110110001111)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0101110110001111) && ({row_reg, col_reg}<16'b0101110110010001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101110110010001) && ({row_reg, col_reg}<16'b0101110110010100)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0101110110010100)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101110110010101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101110110010110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101110110010111) && ({row_reg, col_reg}<16'b0101110110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101110110011010) && ({row_reg, col_reg}<16'b0101110110011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101110110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101110110011101) && ({row_reg, col_reg}<16'b0101110110011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101110110011111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0101110110100000) && ({row_reg, col_reg}<16'b0101110110100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101110110100010) && ({row_reg, col_reg}<16'b0101110110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101110110100110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101110110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101110110101000) && ({row_reg, col_reg}<16'b0101110110101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110110101010) && ({row_reg, col_reg}<16'b0101110110101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101110110101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101110110101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101110110101110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0101110110101111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101110110110000) && ({row_reg, col_reg}<16'b0101110110110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101110110110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101110110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101110110110100) && ({row_reg, col_reg}<16'b0101110110111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110110111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101110110111010) && ({row_reg, col_reg}<16'b0101110110111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110110111100) && ({row_reg, col_reg}<16'b0101110110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101110110111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110111000000) && ({row_reg, col_reg}<16'b0101110111000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110111000010) && ({row_reg, col_reg}<16'b0101110111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110111000110) && ({row_reg, col_reg}<16'b0101110111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110111001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110111001111) && ({row_reg, col_reg}<16'b0101110111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110111010001) && ({row_reg, col_reg}<16'b0101110111101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101110111101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101110111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110111110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101110111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110111110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110111110011) && ({row_reg, col_reg}<16'b0101110111110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110111110111)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0101110111111000) && ({row_reg, col_reg}<16'b0101111000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111000000110) && ({row_reg, col_reg}<16'b0101111000001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101111000001000) && ({row_reg, col_reg}<16'b0101111000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111000001111) && ({row_reg, col_reg}<16'b0101111000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101111000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111000010010) && ({row_reg, col_reg}<16'b0101111000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111000100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111000100110) && ({row_reg, col_reg}<16'b0101111000101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111000101001) && ({row_reg, col_reg}<16'b0101111000101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111000101100) && ({row_reg, col_reg}<16'b0101111000101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101111000101110) && ({row_reg, col_reg}<16'b0101111000110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101111000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111000110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111000110010) && ({row_reg, col_reg}<16'b0101111000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111000110100) && ({row_reg, col_reg}<16'b0101111000110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101111000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101111000110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101111000111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101111000111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101111000111010) && ({row_reg, col_reg}<16'b0101111000111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101111000111100) && ({row_reg, col_reg}<16'b0101111000111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101111000111110) && ({row_reg, col_reg}<16'b0101111001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101111001000001) && ({row_reg, col_reg}<16'b0101111001000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101111001000011) && ({row_reg, col_reg}<16'b0101111001000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101111001000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101111001000111) && ({row_reg, col_reg}<16'b0101111001001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101111001001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101111001001010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101111001001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101111001001100) && ({row_reg, col_reg}<16'b0101111001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111001001111) && ({row_reg, col_reg}<16'b0101111001010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101111001010111) && ({row_reg, col_reg}<16'b0101111001011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111001011010) && ({row_reg, col_reg}<16'b0101111001011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101111001011100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0101111001011101) && ({row_reg, col_reg}<16'b0101111001011111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101111001011111)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0101111001100000)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0101111001100001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101111001100010) && ({row_reg, col_reg}<16'b0101111001100100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101111001100100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101111001100101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0101111001100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101111001100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101111001101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101111001101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111001101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111001101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101111001101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111001101101) && ({row_reg, col_reg}<16'b0101111001110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101111001110000) && ({row_reg, col_reg}<16'b0101111001110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101111001110100) && ({row_reg, col_reg}<16'b0101111001111001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101111001111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101111001111010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0101111001111011) && ({row_reg, col_reg}<16'b0101111001111111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101111001111111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0101111010000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101111010000001) && ({row_reg, col_reg}<16'b0101111010001001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101111010001001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0101111010001010) && ({row_reg, col_reg}<16'b0101111010001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101111010001101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0101111010001110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101111010001111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0101111010010000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101111010010001) && ({row_reg, col_reg}<16'b0101111010010100)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0101111010010100) && ({row_reg, col_reg}<16'b0101111010010110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101111010010110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101111010010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101111010011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101111010011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101111010011010) && ({row_reg, col_reg}<16'b0101111010011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101111010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101111010011101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0101111010011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101111010011111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0101111010100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101111010100001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101111010100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101111010100011) && ({row_reg, col_reg}<16'b0101111010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101111010100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101111010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101111010101000) && ({row_reg, col_reg}<16'b0101111010101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101111010101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101111010101100) && ({row_reg, col_reg}<16'b0101111010101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111010101111) && ({row_reg, col_reg}<16'b0101111010110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101111010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111010110101) && ({row_reg, col_reg}<16'b0101111010110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101111010110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111010111000) && ({row_reg, col_reg}<16'b0101111010111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101111010111010) && ({row_reg, col_reg}<16'b0101111010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101111010111100) && ({row_reg, col_reg}<16'b0101111010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111010111110) && ({row_reg, col_reg}<16'b0101111011000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101111011000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101111011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111011000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101111011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111011000100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111011000101) && ({row_reg, col_reg}<16'b0101111011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111011001001) && ({row_reg, col_reg}<16'b0101111011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101111011001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111011001100) && ({row_reg, col_reg}<16'b0101111011001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111011001111) && ({row_reg, col_reg}<16'b0101111011010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101111011010001) && ({row_reg, col_reg}<16'b0101111011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101111011101101) && ({row_reg, col_reg}<16'b0101111011101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111011101111) && ({row_reg, col_reg}<16'b0101111011110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101111011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111011110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101111011110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111011110100) && ({row_reg, col_reg}<16'b0101111011110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101111011110110) && ({row_reg, col_reg}<16'b0101111011111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111011111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111011111001) && ({row_reg, col_reg}<16'b0101111011111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111011111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101111011111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111011111110)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}>=16'b0101111011111111) && ({row_reg, col_reg}<16'b0101111100000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111100000011) && ({row_reg, col_reg}<16'b0101111100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101111100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111100000110) && ({row_reg, col_reg}<16'b0101111100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101111100001000) && ({row_reg, col_reg}<16'b0101111100001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111100001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111100001111) && ({row_reg, col_reg}<16'b0101111100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111100010010) && ({row_reg, col_reg}<16'b0101111100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101111100100101) && ({row_reg, col_reg}<16'b0101111100101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111100101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111100101010) && ({row_reg, col_reg}<16'b0101111100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101111100101110) && ({row_reg, col_reg}<16'b0101111100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101111100110000) && ({row_reg, col_reg}<16'b0101111100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111100110100) && ({row_reg, col_reg}<16'b0101111100110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101111100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101111100110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101111100111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101111100111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101111100111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101111100111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111100111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101111100111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101111100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111100111111) && ({row_reg, col_reg}<16'b0101111101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101111101000001) && ({row_reg, col_reg}<16'b0101111101000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101111101000100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0101111101000101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101111101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101111101000111) && ({row_reg, col_reg}<16'b0101111101001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101111101001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101111101001010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101111101001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101111101001100) && ({row_reg, col_reg}<16'b0101111101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111101001111) && ({row_reg, col_reg}<16'b0101111101010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101111101010011) && ({row_reg, col_reg}<16'b0101111101010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101111101010111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0101111101011000) && ({row_reg, col_reg}<16'b0101111101011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101111101011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101111101011100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101111101011101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101111101011110) && ({row_reg, col_reg}<16'b0101111101100100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101111101100100) && ({row_reg, col_reg}<16'b0101111101100110)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0101111101100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101111101100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101111101101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101111101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111101101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101111101101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111101101101) && ({row_reg, col_reg}<16'b0101111101110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101111101110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101111101110001) && ({row_reg, col_reg}<16'b0101111101110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101111101110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101111101110100) && ({row_reg, col_reg}<16'b0101111101111100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101111101111100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0101111101111101) && ({row_reg, col_reg}<16'b0101111110001001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101111110001001) && ({row_reg, col_reg}<16'b0101111110001011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101111110001011) && ({row_reg, col_reg}<16'b0101111110001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101111110001101) && ({row_reg, col_reg}<16'b0101111110001111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101111110001111) && ({row_reg, col_reg}<16'b0101111110010001)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101111110010001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101111110010010) && ({row_reg, col_reg}<16'b0101111110010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101111110010101)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0101111110010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101111110010111)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0101111110011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101111110011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101111110011010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101111110011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101111110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101111110011101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0101111110011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101111110011111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0101111110100000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101111110100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101111110100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101111110100011) && ({row_reg, col_reg}<16'b0101111110100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101111110100101) && ({row_reg, col_reg}<16'b0101111110101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101111110101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101111110101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111110101010) && ({row_reg, col_reg}<16'b0101111110110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101111110110000) && ({row_reg, col_reg}<16'b0101111110110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111110110010) && ({row_reg, col_reg}<16'b0101111110110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101111110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111110110101) && ({row_reg, col_reg}<16'b0101111110110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101111110110111) && ({row_reg, col_reg}<16'b0101111110111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101111110111001) && ({row_reg, col_reg}<16'b0101111110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111110111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101111110111111) && ({row_reg, col_reg}<16'b0101111111000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101111111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111111000010) && ({row_reg, col_reg}<16'b0101111111000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111111000101) && ({row_reg, col_reg}<16'b0101111111001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111111001011) && ({row_reg, col_reg}<16'b0101111111001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111111001101) && ({row_reg, col_reg}<16'b0101111111001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111111001111) && ({row_reg, col_reg}<16'b0101111111010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101111111010001) && ({row_reg, col_reg}<16'b0101111111101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111111101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111111101111) && ({row_reg, col_reg}<16'b0101111111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111111110010) && ({row_reg, col_reg}<16'b0101111111110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111111110100) && ({row_reg, col_reg}<16'b0101111111111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111111111100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0101111111111101) && ({row_reg, col_reg}<16'b0110000000000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000000000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110000000000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000000000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110000000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000000000110) && ({row_reg, col_reg}<16'b0110000000001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110000000001000) && ({row_reg, col_reg}<16'b0110000000001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000000001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110000000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000000001101) && ({row_reg, col_reg}<16'b0110000000010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110000000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000000010010) && ({row_reg, col_reg}<16'b0110000000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110000000100101) && ({row_reg, col_reg}<16'b0110000000100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000000100111) && ({row_reg, col_reg}<16'b0110000000101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000000101001) && ({row_reg, col_reg}<16'b0110000000101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110000000101110) && ({row_reg, col_reg}<16'b0110000000110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000000110000) && ({row_reg, col_reg}<16'b0110000000110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000000110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000000110011) && ({row_reg, col_reg}<16'b0110000000110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110000000110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110000000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110000000110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110000000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110000000111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110000000111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110000000111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000000111100) && ({row_reg, col_reg}<16'b0110000000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110000000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000000111111) && ({row_reg, col_reg}<16'b0110000001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110000001000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110000001000010) && ({row_reg, col_reg}<16'b0110000001000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110000001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110000001000110) && ({row_reg, col_reg}<16'b0110000001001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110000001001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110000001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110000001001010) && ({row_reg, col_reg}<16'b0110000001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110000001001100) && ({row_reg, col_reg}<16'b0110000001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110000001001111) && ({row_reg, col_reg}<16'b0110000001010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110000001010011) && ({row_reg, col_reg}<16'b0110000001010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110000001010101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110000001010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110000001010111) && ({row_reg, col_reg}<16'b0110000001011001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110000001011001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110000001011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110000001011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000001011100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110000001011101) && ({row_reg, col_reg}<16'b0110000001011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110000001011111) && ({row_reg, col_reg}<16'b0110000001100001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110000001100001) && ({row_reg, col_reg}<16'b0110000001100011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110000001100011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0110000001100100) && ({row_reg, col_reg}<16'b0110000001100110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110000001100110)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0110000001100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110000001101000)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==16'b0110000001101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110000001101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000001101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110000001101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110000001101101) && ({row_reg, col_reg}<16'b0110000001110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110000001110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110000001110001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110000001110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110000001110011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0110000001110100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110000001110101) && ({row_reg, col_reg}<16'b0110000001111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110000001111010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0110000001111011) && ({row_reg, col_reg}<16'b0110000010000001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110000010000001) && ({row_reg, col_reg}<16'b0110000010001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110000010001000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110000010001001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110000010001010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0110000010001011) && ({row_reg, col_reg}<16'b0110000010001110)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0110000010001110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110000010001111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0110000010010000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110000010010001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110000010010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110000010010011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0110000010010100) && ({row_reg, col_reg}<16'b0110000010011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110000010011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110000010011010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110000010011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110000010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110000010011101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0110000010011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110000010011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000010100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110000010100001) && ({row_reg, col_reg}<16'b0110000010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000010100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110000010100100) && ({row_reg, col_reg}<16'b0110000010101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110000010101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110000010101001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0110000010101010) && ({row_reg, col_reg}<16'b0110000010101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000010101101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110000010101110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110000010101111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110000010110000) && ({row_reg, col_reg}<16'b0110000010110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110000010110010) && ({row_reg, col_reg}<16'b0110000010110100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110000010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110000010110101) && ({row_reg, col_reg}<16'b0110000010110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110000010110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000010111000) && ({row_reg, col_reg}<16'b0110000010111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000010111010) && ({row_reg, col_reg}<16'b0110000010111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110000010111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000010111101) && ({row_reg, col_reg}<16'b0110000011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000011000001) && ({row_reg, col_reg}<16'b0110000011000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000011000011) && ({row_reg, col_reg}<16'b0110000011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000011000110) && ({row_reg, col_reg}<16'b0110000011001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000011001011) && ({row_reg, col_reg}<16'b0110000011001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000011001101) && ({row_reg, col_reg}<16'b0110000011001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000011001111) && ({row_reg, col_reg}<16'b0110000011010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000011010001) && ({row_reg, col_reg}<16'b0110000011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110000011101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000011101111) && ({row_reg, col_reg}<16'b0110000011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000011110001) && ({row_reg, col_reg}<16'b0110000011110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000011110100) && ({row_reg, col_reg}<16'b0110000011110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000011110111)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0110000011111000) && ({row_reg, col_reg}<16'b0110000100000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000100000001) && ({row_reg, col_reg}<16'b0110000100000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110000100000011) && ({row_reg, col_reg}<16'b0110000100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000100000110) && ({row_reg, col_reg}<16'b0110000100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110000100001000) && ({row_reg, col_reg}<16'b0110000100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000100001101) && ({row_reg, col_reg}<16'b0110000100010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110000100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000100010010) && ({row_reg, col_reg}<16'b0110000100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110000100100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000100100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110000100100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000100101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000100101001) && ({row_reg, col_reg}<16'b0110000100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110000100101110) && ({row_reg, col_reg}<16'b0110000100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000100110000) && ({row_reg, col_reg}<16'b0110000100110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000100110010) && ({row_reg, col_reg}<16'b0110000100110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000100110100) && ({row_reg, col_reg}<16'b0110000100110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110000100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110000100110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110000100111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110000100111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110000100111010) && ({row_reg, col_reg}<16'b0110000100111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000100111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110000100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000100111111) && ({row_reg, col_reg}<16'b0110000101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000101000001) && ({row_reg, col_reg}<16'b0110000101000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110000101000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110000101000100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0110000101000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110000101000110) && ({row_reg, col_reg}<16'b0110000101001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110000101001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110000101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110000101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110000101001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110000101001101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110000101001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110000101001111) && ({row_reg, col_reg}<16'b0110000101010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000101010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110000101010011) && ({row_reg, col_reg}<16'b0110000101010111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110000101010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110000101011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000101011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110000101011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110000101011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000101011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110000101011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110000101011110) && ({row_reg, col_reg}<16'b0110000101100011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110000101100011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110000101100100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110000101100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110000101100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110000101100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110000101101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110000101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110000101101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110000101101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110000101101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110000101101101) && ({row_reg, col_reg}<16'b0110000101110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110000101110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110000101110001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110000101110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110000101110011) && ({row_reg, col_reg}<16'b0110000101110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0110000101110101) && ({row_reg, col_reg}<16'b0110000101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000101111011) && ({row_reg, col_reg}<16'b0110000110000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110000110000001) && ({row_reg, col_reg}<16'b0110000110000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110000110000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110000110000101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110000110000110) && ({row_reg, col_reg}<16'b0110000110001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110000110001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110000110001001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0110000110001010) && ({row_reg, col_reg}<16'b0110000110001100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0110000110001100) && ({row_reg, col_reg}<16'b0110000110001111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0110000110001111) && ({row_reg, col_reg}<16'b0110000110010010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0110000110010010) && ({row_reg, col_reg}<16'b0110000110010101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110000110010101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0110000110010110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110000110010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110000110011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000110011001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110000110011010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110000110011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110000110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110000110011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000110011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110000110011111) && ({row_reg, col_reg}<16'b0110000110100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110000110100011) && ({row_reg, col_reg}<16'b0110000110100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110000110100101) && ({row_reg, col_reg}<16'b0110000110100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110000110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110000110101000) && ({row_reg, col_reg}<16'b0110000110101010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110000110101010) && ({row_reg, col_reg}<16'b0110000110101110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110000110101110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110000110101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110000110110000) && ({row_reg, col_reg}<16'b0110000110110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110000110110010) && ({row_reg, col_reg}<16'b0110000110110100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110000110110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110000110110101) && ({row_reg, col_reg}<16'b0110000110110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110000110110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110000110111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000110111001) && ({row_reg, col_reg}<16'b0110000110111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110000110111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000110111101) && ({row_reg, col_reg}<16'b0110000110111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110000110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110000111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000111000001) && ({row_reg, col_reg}<16'b0110000111000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000111000011) && ({row_reg, col_reg}<16'b0110000111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000111000110) && ({row_reg, col_reg}<16'b0110000111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000111001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110000111001001) && ({row_reg, col_reg}<16'b0110000111001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000111001011) && ({row_reg, col_reg}<16'b0110000111001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110000111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000111001111) && ({row_reg, col_reg}<16'b0110000111010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000111010001) && ({row_reg, col_reg}<16'b0110000111101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110000111101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000111101111) && ({row_reg, col_reg}<16'b0110000111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000111110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110000111110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110000111110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000111110100) && ({row_reg, col_reg}<16'b0110000111111001)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0110000111111001) && ({row_reg, col_reg}<16'b0110001000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001000000000) && ({row_reg, col_reg}<16'b0110001000001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110001000001000) && ({row_reg, col_reg}<16'b0110001000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001000001101) && ({row_reg, col_reg}<16'b0110001000010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110001000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001000010010) && ({row_reg, col_reg}<16'b0110001000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110001000100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001000100110) && ({row_reg, col_reg}<16'b0110001000101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110001000101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001000101001) && ({row_reg, col_reg}<16'b0110001000101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110001000101110) && ({row_reg, col_reg}<16'b0110001000110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110001000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001000110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001000110010) && ({row_reg, col_reg}<16'b0110001000110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001000110100) && ({row_reg, col_reg}<16'b0110001000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110001000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001000110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110001000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001000111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110001000111010) && ({row_reg, col_reg}<16'b0110001000111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001000111111) && ({row_reg, col_reg}<16'b0110001001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001001000001) && ({row_reg, col_reg}<16'b0110001001000101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110001001000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001001000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110001001000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001001001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110001001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110001001001100) && ({row_reg, col_reg}<16'b0110001001001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110001001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110001001001111) && ({row_reg, col_reg}<16'b0110001001010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110001001010010) && ({row_reg, col_reg}<16'b0110001001010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001001010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110001001010101) && ({row_reg, col_reg}<16'b0110001001010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001001010111) && ({row_reg, col_reg}<16'b0110001001011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001001011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110001001011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001001011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001001011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001001011110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0110001001011111) && ({row_reg, col_reg}<16'b0110001001100001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110001001100001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0110001001100010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110001001100011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110001001100100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110001001100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110001001100110) && ({row_reg, col_reg}<16'b0110001001101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001001101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001001101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110001001101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001001101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110001001101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110001001101101) && ({row_reg, col_reg}<16'b0110001001110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110001001110000) && ({row_reg, col_reg}<16'b0110001001110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110001001110011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110001001110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0110001001110101) && ({row_reg, col_reg}<16'b0110001001111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001001111101) && ({row_reg, col_reg}<16'b0110001001111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0110001001111111) && ({row_reg, col_reg}<16'b0110001010000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110001010000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001010000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110001010000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110001010000110) && ({row_reg, col_reg}<16'b0110001010001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110001010001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110001010001001)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0110001010001010)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0110001010001011) && ({row_reg, col_reg}<16'b0110001010001111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0110001010001111) && ({row_reg, col_reg}<16'b0110001010010001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110001010010001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110001010010010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110001010010011)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0110001010010100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110001010010101)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0110001010010110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110001010010111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110001010011000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110001010011001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110001010011010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110001010011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110001010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110001010011101) && ({row_reg, col_reg}<16'b0110001010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110001010100011) && ({row_reg, col_reg}<16'b0110001010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110001010100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001010100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110001010101000) && ({row_reg, col_reg}<16'b0110001010101010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110001010101010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0110001010101011) && ({row_reg, col_reg}<16'b0110001010101110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110001010101110) && ({row_reg, col_reg}<16'b0110001010110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001010110000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110001010110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001010110010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0110001010110011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110001010110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110001010110101) && ({row_reg, col_reg}<16'b0110001010110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110001010110111) && ({row_reg, col_reg}<16'b0110001010111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001010111001) && ({row_reg, col_reg}<16'b0110001010111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110001010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001010111110) && ({row_reg, col_reg}<16'b0110001011000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110001011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001011000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001011000010) && ({row_reg, col_reg}<16'b0110001011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110001011000100) && ({row_reg, col_reg}<16'b0110001011000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001011000111) && ({row_reg, col_reg}<16'b0110001011001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110001011001001) && ({row_reg, col_reg}<16'b0110001011001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110001011001100) && ({row_reg, col_reg}<16'b0110001011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110001011001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110001011001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110001011010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001011010001) && ({row_reg, col_reg}<16'b0110001011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110001011101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001011101111) && ({row_reg, col_reg}<16'b0110001011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001011110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001011110010) && ({row_reg, col_reg}<16'b0110001011110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110001011110100) && ({row_reg, col_reg}<16'b0110001011111011)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0110001011111011) && ({row_reg, col_reg}<16'b0110001100000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001100000001) && ({row_reg, col_reg}<16'b0110001100000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110001100000011) && ({row_reg, col_reg}<16'b0110001100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001100000101) && ({row_reg, col_reg}<16'b0110001100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110001100001000) && ({row_reg, col_reg}<16'b0110001100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001100001101) && ({row_reg, col_reg}<16'b0110001100010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110001100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001100010010) && ({row_reg, col_reg}<16'b0110001100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110001100100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001100100110) && ({row_reg, col_reg}<16'b0110001100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110001100101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001100101001) && ({row_reg, col_reg}<16'b0110001100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110001100101110) && ({row_reg, col_reg}<16'b0110001100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001100110000) && ({row_reg, col_reg}<16'b0110001100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001100110100) && ({row_reg, col_reg}<16'b0110001100110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110001100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001100110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110001100111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001100111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110001100111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001100111011) && ({row_reg, col_reg}<16'b0110001101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001101000100) && ({row_reg, col_reg}<16'b0110001101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001101000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110001101000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001101001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110001101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110001101001011) && ({row_reg, col_reg}<16'b0110001101001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001101001101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0110001101001110) && ({row_reg, col_reg}<16'b0110001101010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001101010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001101010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001101010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110001101010101) && ({row_reg, col_reg}<16'b0110001101010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110001101010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001101011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110001101011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001101011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110001101011011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0110001101011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001101011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110001101011110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110001101011111)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}>=16'b0110001101100000) && ({row_reg, col_reg}<16'b0110001101100010)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0110001101100010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110001101100011)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0110001101100100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110001101100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110001101100110)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0110001101100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110001101101000) && ({row_reg, col_reg}<16'b0110001101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001101101011) && ({row_reg, col_reg}<16'b0110001101101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110001101101101) && ({row_reg, col_reg}<16'b0110001101110001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110001101110001) && ({row_reg, col_reg}<16'b0110001101110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0110001101110011) && ({row_reg, col_reg}<16'b0110001101110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110001101110111)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}>=16'b0110001101111000) && ({row_reg, col_reg}<16'b0110001101111011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110001101111011)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}>=16'b0110001101111100) && ({row_reg, col_reg}<16'b0110001110000010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110001110000010)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}>=16'b0110001110000011) && ({row_reg, col_reg}<16'b0110001110000111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110001110000111)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}>=16'b0110001110001000) && ({row_reg, col_reg}<16'b0110001110001010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110001110001010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110001110001011)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0110001110001100) && ({row_reg, col_reg}<16'b0110001110001110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110001110001110)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0110001110001111) && ({row_reg, col_reg}<16'b0110001110010001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0110001110010001) && ({row_reg, col_reg}<16'b0110001110010110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110001110010110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110001110010111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0110001110011000) && ({row_reg, col_reg}<16'b0110001110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001110011010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110001110011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110001110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110001110011101) && ({row_reg, col_reg}<16'b0110001110100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001110100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110001110100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110001110100011) && ({row_reg, col_reg}<16'b0110001110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110001110100110) && ({row_reg, col_reg}<16'b0110001110101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110001110101000) && ({row_reg, col_reg}<16'b0110001110101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110001110101011) && ({row_reg, col_reg}<16'b0110001110101110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001110101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001110101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110001110110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110001110110001) && ({row_reg, col_reg}<16'b0110001110110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110001110110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110001110110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110001110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001110111001) && ({row_reg, col_reg}<16'b0110001110111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110001110111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110001110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001110111110) && ({row_reg, col_reg}<16'b0110001111000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110001111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001111000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001111000010) && ({row_reg, col_reg}<16'b0110001111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110001111000100) && ({row_reg, col_reg}<16'b0110001111001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001111001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001111001100) && ({row_reg, col_reg}<16'b0110001111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001111001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001111001111) && ({row_reg, col_reg}<16'b0110001111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001111010001) && ({row_reg, col_reg}<16'b0110001111101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110001111101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001111101111) && ({row_reg, col_reg}<16'b0110001111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001111110010) && ({row_reg, col_reg}<16'b0110001111110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001111110110) && ({row_reg, col_reg}<16'b0110001111111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001111111011) && ({row_reg, col_reg}<16'b0110001111111110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0110001111111110) && ({row_reg, col_reg}<16'b0110010000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110010000000000) && ({row_reg, col_reg}<16'b0110010000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010000000110) && ({row_reg, col_reg}<16'b0110010000001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110010000001000) && ({row_reg, col_reg}<16'b0110010000001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010000001110) && ({row_reg, col_reg}<16'b0110010000010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110010000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010000010010) && ({row_reg, col_reg}<16'b0110010000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110010000100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010000100110) && ({row_reg, col_reg}<16'b0110010000101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110010000101001) && ({row_reg, col_reg}<16'b0110010000101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110010000101110) && ({row_reg, col_reg}<16'b0110010000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010000110001) && ({row_reg, col_reg}<16'b0110010000110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110010000110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010000110100) && ({row_reg, col_reg}<16'b0110010000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110010000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110010000110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110010000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110010000111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110010000111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010000111011) && ({row_reg, col_reg}<16'b0110010001000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010001000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110010001000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110010001000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110010001000111) && ({row_reg, col_reg}<16'b0110010001001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110010001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110010001001010) && ({row_reg, col_reg}<16'b0110010001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110010001001100) && ({row_reg, col_reg}<16'b0110010001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110010001001111) && ({row_reg, col_reg}<16'b0110010001010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110010001010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110010001010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110010001010101) && ({row_reg, col_reg}<16'b0110010001010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010001010111) && ({row_reg, col_reg}<16'b0110010001011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110010001011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010001011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110010001011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110010001011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110010001011110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110010001011111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110010001100000)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0110010001100001) && ({row_reg, col_reg}<16'b0110010001100011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110010001100011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110010001100100)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0110010001100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110010001100110) && ({row_reg, col_reg}<16'b0110010001101000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0110010001101000) && ({row_reg, col_reg}<16'b0110010001101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110010001101011) && ({row_reg, col_reg}<16'b0110010001110111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0110010001110111) && ({row_reg, col_reg}<16'b0110010001111110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110010001111110) && ({row_reg, col_reg}<16'b0110010010000001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0110010010000001) && ({row_reg, col_reg}<16'b0110010010000011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0110010010000011) && ({row_reg, col_reg}<16'b0110010010000110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110010010000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110010010000111)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0110010010001000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110010010001001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110010010001010)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0110010010001011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110010010001100)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}>=16'b0110010010001101) && ({row_reg, col_reg}<16'b0110010010001111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110010010001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110010010010000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110010010010001)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}>=16'b0110010010010010) && ({row_reg, col_reg}<16'b0110010010010111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110010010010111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0110010010011000) && ({row_reg, col_reg}<16'b0110010010011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110010010011100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110010010011101) && ({row_reg, col_reg}<16'b0110010010100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110010010100000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110010010100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110010010100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110010010100011) && ({row_reg, col_reg}<16'b0110010010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110010010100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110010010100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110010010101000) && ({row_reg, col_reg}<16'b0110010010101010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0110010010101010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110010010101011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0110010010101100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110010010101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110010010101110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110010010101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110010010110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110010010110001) && ({row_reg, col_reg}<16'b0110010010110011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110010010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110010010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110010010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110010010110110) && ({row_reg, col_reg}<16'b0110010010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110010010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010010111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010010111010) && ({row_reg, col_reg}<16'b0110010010111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110010010111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110010010111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010010111110) && ({row_reg, col_reg}<16'b0110010011000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110010011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010011000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010011000010) && ({row_reg, col_reg}<16'b0110010011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110010011000100) && ({row_reg, col_reg}<16'b0110010011001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110010011001100) && ({row_reg, col_reg}<16'b0110010011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010011001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110010011001111) && ({row_reg, col_reg}<16'b0110010011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010011010001) && ({row_reg, col_reg}<16'b0110010011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110010011101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110010011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010011110010) && ({row_reg, col_reg}<16'b0110010011110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110010011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110010011110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010011110111) && ({row_reg, col_reg}<16'b0110010011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010011111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010011111010) && ({row_reg, col_reg}<16'b0110010011111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110010011111100) && ({row_reg, col_reg}<16'b0110010011111110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0110010011111110) && ({row_reg, col_reg}<16'b0110010100000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110010100000001) && ({row_reg, col_reg}<16'b0110010100000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010100000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110010100000101) && ({row_reg, col_reg}<16'b0110010100000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010100000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110010100001000) && ({row_reg, col_reg}<16'b0110010100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010100010010) && ({row_reg, col_reg}<16'b0110010100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110010100100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010100100110) && ({row_reg, col_reg}<16'b0110010100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110010100101001) && ({row_reg, col_reg}<16'b0110010100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110010100101110) && ({row_reg, col_reg}<16'b0110010100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010100110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110010100110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110010100110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110010100110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010100110100) && ({row_reg, col_reg}<16'b0110010100110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110010100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110010100110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110010100111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110010100111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110010100111010) && ({row_reg, col_reg}<16'b0110010100111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010100111100) && ({row_reg, col_reg}<16'b0110010101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010101000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110010101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110010101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110010101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110010101000111) && ({row_reg, col_reg}<16'b0110010101001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110010101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110010101001010) && ({row_reg, col_reg}<16'b0110010101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110010101001100) && ({row_reg, col_reg}<16'b0110010101001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110010101001110) && ({row_reg, col_reg}<16'b0110010101010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110010101010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110010101010011) && ({row_reg, col_reg}<16'b0110010101010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110010101010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010101010110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010101010111) && ({row_reg, col_reg}<16'b0110010101011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110010101011010)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==16'b0110010101011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010101011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110010101011101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0110010101011110)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0110010101011111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110010101100000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0110010101100001) && ({row_reg, col_reg}<16'b0110010101100011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110010101100011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0110010101100100) && ({row_reg, col_reg}<16'b0110010101101000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110010101101000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0110010101101001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110010101101010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0110010101101011) && ({row_reg, col_reg}<16'b0110010101110100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110010101110100)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0110010101110101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110010101110110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0110010101110111) && ({row_reg, col_reg}<16'b0110010101111110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110010101111110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110010101111111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110010110000000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0110010110000001) && ({row_reg, col_reg}<16'b0110010110000011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110010110000011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110010110000100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110010110000101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0110010110000110) && ({row_reg, col_reg}<16'b0110010110001001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110010110001001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110010110001010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110010110001011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110010110001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110010110001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110010110001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110010110001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110010110010000) && ({row_reg, col_reg}<16'b0110010110011010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110010110011010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110010110011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110010110011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110010110011101) && ({row_reg, col_reg}<16'b0110010110100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110010110100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110010110100001) && ({row_reg, col_reg}<16'b0110010110100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110010110100011) && ({row_reg, col_reg}<16'b0110010110100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110010110100111) && ({row_reg, col_reg}<16'b0110010110101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110010110101011) && ({row_reg, col_reg}<16'b0110010110101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110010110101101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110010110101110) && ({row_reg, col_reg}<16'b0110010110110001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110010110110001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110010110110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110010110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110010110110100) && ({row_reg, col_reg}<16'b0110010110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110010110111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110010110111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010110111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110010110111011) && ({row_reg, col_reg}<16'b0110010110111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110010110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010110111110) && ({row_reg, col_reg}<16'b0110010111000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110010111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010111000010) && ({row_reg, col_reg}<16'b0110010111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110010111000100) && ({row_reg, col_reg}<16'b0110010111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010111000111) && ({row_reg, col_reg}<16'b0110010111001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010111001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010111001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110010111001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110010111001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110010111001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010111001111) && ({row_reg, col_reg}<16'b0110010111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010111010001) && ({row_reg, col_reg}<16'b0110010111101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110010111101111) && ({row_reg, col_reg}<16'b0110010111110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010111110010) && ({row_reg, col_reg}<16'b0110010111110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110010111110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010111110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110010111111000) && ({row_reg, col_reg}<16'b0110010111111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010111111010) && ({row_reg, col_reg}<16'b0110010111111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010111111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010111111101)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}>=16'b0110010111111110) && ({row_reg, col_reg}<16'b0110011000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011000000000) && ({row_reg, col_reg}<16'b0110011000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011000010011) && ({row_reg, col_reg}<16'b0110011000100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110011000100100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110011000100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011000100110) && ({row_reg, col_reg}<16'b0110011000101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110011000101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011000101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011000101010) && ({row_reg, col_reg}<16'b0110011000101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110011000101110) && ({row_reg, col_reg}<16'b0110011000110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110011000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011000110001) && ({row_reg, col_reg}<16'b0110011000110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110011000110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011000110100) && ({row_reg, col_reg}<16'b0110011000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110011000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110011000110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110011000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110011000111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110011000111010) && ({row_reg, col_reg}<16'b0110011000111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011000111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110011000111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110011000111110) && ({row_reg, col_reg}<16'b0110011001000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011001000010) && ({row_reg, col_reg}<16'b0110011001000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0110011001000100) && ({row_reg, col_reg}<16'b0110011001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110011001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110011001000111) && ({row_reg, col_reg}<16'b0110011001001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110011001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110011001001010) && ({row_reg, col_reg}<16'b0110011001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110011001001100) && ({row_reg, col_reg}<16'b0110011001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110011001001110) && ({row_reg, col_reg}<16'b0110011001010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110011001010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110011001010011) && ({row_reg, col_reg}<16'b0110011001010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110011001010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011001010110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011001010111) && ({row_reg, col_reg}<16'b0110011001011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110011001011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110011001011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110011001011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110011001011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011001011110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110011001011111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110011001100000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0110011001100001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110011001100010)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0110011001100011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0110011001100100) && ({row_reg, col_reg}<16'b0110011001100110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0110011001100110) && ({row_reg, col_reg}<16'b0110011001101000)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0110011001101000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110011001101001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0110011001101010)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0110011001101011) && ({row_reg, col_reg}<16'b0110011001101110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110011001101110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0110011001101111) && ({row_reg, col_reg}<16'b0110011001110100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110011001110100)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0110011001110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110011001110110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110011001110111)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}>=16'b0110011001111000) && ({row_reg, col_reg}<16'b0110011001111100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110011001111100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0110011001111101) && ({row_reg, col_reg}<16'b0110011001111111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110011001111111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110011010000000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0110011010000001) && ({row_reg, col_reg}<16'b0110011010000100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0110011010000100) && ({row_reg, col_reg}<16'b0110011010001000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110011010001000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110011010001001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110011010001010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110011010001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110011010001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110011010001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011010001110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110011010001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110011010010000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0110011010010001) && ({row_reg, col_reg}<16'b0110011010010011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110011010010011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0110011010010100) && ({row_reg, col_reg}<16'b0110011010011001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110011010011001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110011010011010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110011010011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011010011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110011010011101) && ({row_reg, col_reg}<16'b0110011010100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110011010100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110011010100001) && ({row_reg, col_reg}<16'b0110011010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110011010100011) && ({row_reg, col_reg}<16'b0110011010100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110011010100111) && ({row_reg, col_reg}<16'b0110011010101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110011010101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110011010101100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0110011010101101) && ({row_reg, col_reg}<16'b0110011010110000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110011010110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110011010110001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110011010110010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110011010110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011010110100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0110011010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110011010110110) && ({row_reg, col_reg}<16'b0110011010111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110011010111000) && ({row_reg, col_reg}<16'b0110011010111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011010111010) && ({row_reg, col_reg}<16'b0110011010111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011010111100) && ({row_reg, col_reg}<16'b0110011010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011010111110) && ({row_reg, col_reg}<16'b0110011011000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110011011000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110011011000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011011000010) && ({row_reg, col_reg}<16'b0110011011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110011011000100) && ({row_reg, col_reg}<16'b0110011011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011011000110) && ({row_reg, col_reg}<16'b0110011011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011011001000) && ({row_reg, col_reg}<16'b0110011011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011011001010) && ({row_reg, col_reg}<16'b0110011011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011011010001) && ({row_reg, col_reg}<16'b0110011011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110011011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110011011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011011110010) && ({row_reg, col_reg}<16'b0110011011110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110011011110111)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0110011011111000) && ({row_reg, col_reg}<16'b0110011100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011100000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110011100000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011100000011) && ({row_reg, col_reg}<16'b0110011100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011100010011) && ({row_reg, col_reg}<16'b0110011100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110011100100101) && ({row_reg, col_reg}<16'b0110011100100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011100100111) && ({row_reg, col_reg}<16'b0110011100101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011100101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011100101010) && ({row_reg, col_reg}<16'b0110011100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110011100101110) && ({row_reg, col_reg}<16'b0110011100110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011100110001) && ({row_reg, col_reg}<16'b0110011100110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110011100110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011100110100) && ({row_reg, col_reg}<16'b0110011100110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110011100110110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0110011100110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110011100111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110011100111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110011100111010) && ({row_reg, col_reg}<16'b0110011100111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011100111100) && ({row_reg, col_reg}<16'b0110011100111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110011100111110) && ({row_reg, col_reg}<16'b0110011101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110011101000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110011101000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110011101000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110011101000100) && ({row_reg, col_reg}<16'b0110011101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110011101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110011101000111) && ({row_reg, col_reg}<16'b0110011101001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110011101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110011101001010) && ({row_reg, col_reg}<16'b0110011101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110011101001100) && ({row_reg, col_reg}<16'b0110011101001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110011101001110) && ({row_reg, col_reg}<16'b0110011101010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110011101010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110011101010011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110011101010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110011101010101) && ({row_reg, col_reg}<16'b0110011101010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011101010111) && ({row_reg, col_reg}<16'b0110011101011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110011101011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011101011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110011101011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110011101011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110011101011110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110011101011111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110011101100000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0110011101100001) && ({row_reg, col_reg}<16'b0110011101100011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110011101100011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0110011101100100) && ({row_reg, col_reg}<16'b0110011101101000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110011101101000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0110011101101001) && ({row_reg, col_reg}<16'b0110011101101011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110011101101011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0110011101101100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110011101101101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110011101101110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110011101101111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110011101110000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0110011101110001) && ({row_reg, col_reg}<16'b0110011101110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110011101110011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110011101110100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110011101110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110011101110110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0110011101110111) && ({row_reg, col_reg}<16'b0110011101111011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110011101111011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110011101111100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110011101111101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110011101111110)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0110011101111111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110011110000000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0110011110000001) && ({row_reg, col_reg}<16'b0110011110000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110011110000100) && ({row_reg, col_reg}<16'b0110011110000111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110011110000111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110011110001000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110011110001001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110011110001010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110011110001011) && ({row_reg, col_reg}<16'b0110011110001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110011110001101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110011110001110) && ({row_reg, col_reg}<16'b0110011110010000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110011110010000) && ({row_reg, col_reg}<16'b0110011110010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011110010011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110011110010100) && ({row_reg, col_reg}<16'b0110011110011000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110011110011000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110011110011001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110011110011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110011110011011) && ({row_reg, col_reg}<16'b0110011110011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110011110011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110011110100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110011110100001) && ({row_reg, col_reg}<16'b0110011110100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110011110100011) && ({row_reg, col_reg}<16'b0110011110100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110011110100111) && ({row_reg, col_reg}<16'b0110011110101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110011110101001) && ({row_reg, col_reg}<16'b0110011110101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110011110101011) && ({row_reg, col_reg}<16'b0110011110101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110011110101101) && ({row_reg, col_reg}<16'b0110011110110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011110110010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110011110110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011110110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0110011110110101) && ({row_reg, col_reg}<16'b0110011110110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011110110111) && ({row_reg, col_reg}<16'b0110011110111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110011110111001) && ({row_reg, col_reg}<16'b0110011110111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011110111100) && ({row_reg, col_reg}<16'b0110011110111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011110111110) && ({row_reg, col_reg}<16'b0110011111000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110011111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011111000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011111000010) && ({row_reg, col_reg}<16'b0110011111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110011111000100) && ({row_reg, col_reg}<16'b0110011111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110011111000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011111000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110011111001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110011111001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011111001010) && ({row_reg, col_reg}<16'b0110011111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011111010001) && ({row_reg, col_reg}<16'b0110011111110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110011111110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011111111000) && ({row_reg, col_reg}<16'b0110011111111111)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}==16'b0110011111111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110100000000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110100000000001) && ({row_reg, col_reg}<16'b0110100000001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100000001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100000001111) && ({row_reg, col_reg}<16'b0110100000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100000010010) && ({row_reg, col_reg}<16'b0110100000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110100000100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100000100110) && ({row_reg, col_reg}<16'b0110100000101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100000101000) && ({row_reg, col_reg}<16'b0110100000101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100000101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100000101011) && ({row_reg, col_reg}<16'b0110100000101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110100000101101) && ({row_reg, col_reg}<16'b0110100000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100000110001) && ({row_reg, col_reg}<16'b0110100000110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110100000110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100000110100) && ({row_reg, col_reg}<16'b0110100000110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110100000110111) && ({row_reg, col_reg}<16'b0110100000111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110100000111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110100000111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110100000111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100000111100) && ({row_reg, col_reg}<16'b0110100000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110100000111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100000111111) && ({row_reg, col_reg}<16'b0110100001000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110100001000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110100001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110100001000110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0110100001000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110100001001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110100001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110100001001010) && ({row_reg, col_reg}<16'b0110100001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110100001001100) && ({row_reg, col_reg}<16'b0110100001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110100001001111) && ({row_reg, col_reg}<16'b0110100001010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110100001010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110100001010100) && ({row_reg, col_reg}<16'b0110100001010110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110100001010110) && ({row_reg, col_reg}<16'b0110100001011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100001011000) && ({row_reg, col_reg}<16'b0110100001011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100001011010) && ({row_reg, col_reg}<16'b0110100001011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110100001011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110100001011101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0110100001011110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110100001011111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0110100001100000) && ({row_reg, col_reg}<16'b0110100001100010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110100001100010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110100001100011) && ({row_reg, col_reg}<16'b0110100001100101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110100001100101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0110100001100110) && ({row_reg, col_reg}<16'b0110100001101000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110100001101000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0110100001101001) && ({row_reg, col_reg}<16'b0110100001101011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110100001101011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0110100001101100) && ({row_reg, col_reg}<16'b0110100001101110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110100001101110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0110100001101111) && ({row_reg, col_reg}<16'b0110100001110001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0110100001110001) && ({row_reg, col_reg}<16'b0110100001110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110100001110011) && ({row_reg, col_reg}<16'b0110100001110101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110100001110101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0110100001110110) && ({row_reg, col_reg}<16'b0110100001111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110100001111000) && ({row_reg, col_reg}<16'b0110100001111010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110100001111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110100001111011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0110100001111100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110100001111101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0110100001111110) && ({row_reg, col_reg}<16'b0110100010000000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110100010000000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0110100010000001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110100010000010)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0110100010000011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110100010000100)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0110100010000101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110100010000110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0110100010000111) && ({row_reg, col_reg}<16'b0110100010001001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110100010001001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110100010001010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110100010001011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0110100010001100) && ({row_reg, col_reg}<16'b0110100010001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110100010001110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110100010001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110100010010000) && ({row_reg, col_reg}<16'b0110100010010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110100010010010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110100010010011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110100010010100) && ({row_reg, col_reg}<16'b0110100010011000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110100010011000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110100010011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110100010011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110100010011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100010011100) && ({row_reg, col_reg}<16'b0110100010011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110100010011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110100010011111) && ({row_reg, col_reg}<16'b0110100010100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110100010100010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0110100010100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110100010100100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0110100010100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110100010100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0110100010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110100010101000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0110100010101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110100010101010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0110100010101011) && ({row_reg, col_reg}<16'b0110100010101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110100010101101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0110100010101110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110100010101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110100010110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110100010110001) && ({row_reg, col_reg}<16'b0110100010110011)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0110100010110011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110100010110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110100010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110100010110110) && ({row_reg, col_reg}<16'b0110100010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110100010111000) && ({row_reg, col_reg}<16'b0110100010111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110100010111010) && ({row_reg, col_reg}<16'b0110100011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110100011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100011000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100011000010) && ({row_reg, col_reg}<16'b0110100011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110100011000100) && ({row_reg, col_reg}<16'b0110100011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110100011000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100011000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110100011001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110100011001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100011001010) && ({row_reg, col_reg}<16'b0110100011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100011001111) && ({row_reg, col_reg}<16'b0110100011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100011010001) && ({row_reg, col_reg}<16'b0110100011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110100011101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100011101110) && ({row_reg, col_reg}<16'b0110100011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110100011110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100011110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100011111000) && ({row_reg, col_reg}<16'b0110100011111111)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}==16'b0110100011111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110100100000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110100100000001) && ({row_reg, col_reg}<16'b0110100100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100100000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110100100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100100000111) && ({row_reg, col_reg}<16'b0110100100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100100001001) && ({row_reg, col_reg}<16'b0110100100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100100001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110100100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110100100001111) && ({row_reg, col_reg}<16'b0110100100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100100010010) && ({row_reg, col_reg}<16'b0110100100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110100100100110) && ({row_reg, col_reg}<16'b0110100100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100100101001) && ({row_reg, col_reg}<16'b0110100100110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100100110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110100100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110100100110011) && ({row_reg, col_reg}<16'b0110100100110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100100110110) && ({row_reg, col_reg}<16'b0110100100111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110100100111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110100100111010) && ({row_reg, col_reg}<16'b0110100100111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110100100111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110100100111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110100100111110) && ({row_reg, col_reg}<16'b0110100101000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100101000000) && ({row_reg, col_reg}<16'b0110100101000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110100101000100) && ({row_reg, col_reg}<16'b0110100101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110100101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110100101000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100101001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110100101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110100101001010) && ({row_reg, col_reg}<16'b0110100101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110100101001100) && ({row_reg, col_reg}<16'b0110100101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110100101001111) && ({row_reg, col_reg}<16'b0110100101010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110100101010011) && ({row_reg, col_reg}<16'b0110100101010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110100101010101) && ({row_reg, col_reg}<16'b0110100101010111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110100101010111) && ({row_reg, col_reg}<16'b0110100101011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100101011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110100101011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110100101011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110100101011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110100101011110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110100101011111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0110100101100000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110100101100001)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0110100101100010)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0110100101100011) && ({row_reg, col_reg}<16'b0110100101100101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0110100101100101) && ({row_reg, col_reg}<16'b0110100101101000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110100101101000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0110100101101001) && ({row_reg, col_reg}<16'b0110100101101100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110100101101100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110100101101101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0110100101101110) && ({row_reg, col_reg}<16'b0110100101110001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0110100101110001) && ({row_reg, col_reg}<16'b0110100101110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110100101110011) && ({row_reg, col_reg}<16'b0110100101110110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0110100101110110) && ({row_reg, col_reg}<16'b0110100101111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110100101111000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110100101111001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110100101111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110100101111011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0110100101111100) && ({row_reg, col_reg}<16'b0110100110000000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110100110000000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110100110000001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110100110000010) && ({row_reg, col_reg}<16'b0110100110000100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110100110000100)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0110100110000101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110100110000110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110100110000111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110100110001000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0110100110001001) && ({row_reg, col_reg}<16'b0110100110001011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110100110001011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110100110001100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110100110001101) && ({row_reg, col_reg}<16'b0110100110001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110100110001111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110100110010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110100110010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110100110010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110100110010011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110100110010100) && ({row_reg, col_reg}<16'b0110100110011000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110100110011000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110100110011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110100110011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110100110011011) && ({row_reg, col_reg}<16'b0110100110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110100110011101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==16'b0110100110011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110100110011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110100110100000) && ({row_reg, col_reg}<16'b0110100110100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110100110100010) && ({row_reg, col_reg}<16'b0110100110100100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110100110100100)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0110100110100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110100110100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0110100110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110100110101000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0110100110101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110100110101010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0110100110101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110100110101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110100110101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110100110101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110100110101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110100110110000) && ({row_reg, col_reg}<16'b0110100110110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110100110110010)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0110100110110011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110100110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110100110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110100110110110) && ({row_reg, col_reg}<16'b0110100110111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110100110111011) && ({row_reg, col_reg}<16'b0110100110111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110100110111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110100110111111) && ({row_reg, col_reg}<16'b0110100111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100111000001) && ({row_reg, col_reg}<16'b0110100111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110100111000100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100111000101) && ({row_reg, col_reg}<16'b0110100111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100111001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100111001111) && ({row_reg, col_reg}<16'b0110100111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100111010001) && ({row_reg, col_reg}<16'b0110100111101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110100111101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100111101110) && ({row_reg, col_reg}<16'b0110100111110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110100111110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100111110111) && ({row_reg, col_reg}<16'b0110100111111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100111111001) && ({row_reg, col_reg}<16'b0110100111111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100111111110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0110100111111111) && ({row_reg, col_reg}<16'b0110101000000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101000000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110101000000010) && ({row_reg, col_reg}<16'b0110101000000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101000000111) && ({row_reg, col_reg}<16'b0110101000001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110101000001010) && ({row_reg, col_reg}<16'b0110101000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101000001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110101000001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110101000001111) && ({row_reg, col_reg}<16'b0110101000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110101000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101000010010) && ({row_reg, col_reg}<16'b0110101000100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110101000100110) && ({row_reg, col_reg}<16'b0110101000101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110101000101001) && ({row_reg, col_reg}<16'b0110101000101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101000101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110101000101100) && ({row_reg, col_reg}<16'b0110101000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101000110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110101000110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110101000110011) && ({row_reg, col_reg}<16'b0110101000110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110101000110111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0110101000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110101000111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110101000111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110101000111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110101000111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110101000111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110101000111110) && ({row_reg, col_reg}<16'b0110101001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110101001000001) && ({row_reg, col_reg}<16'b0110101001000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110101001000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110101001000100) && ({row_reg, col_reg}<16'b0110101001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101001000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110101001000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110101001001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110101001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110101001001010) && ({row_reg, col_reg}<16'b0110101001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110101001001100) && ({row_reg, col_reg}<16'b0110101001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110101001001111) && ({row_reg, col_reg}<16'b0110101001010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101001010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110101001010110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110101001010111) && ({row_reg, col_reg}<16'b0110101001011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101001011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110101001011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110101001011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110101001011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110101001011110)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}>=16'b0110101001011111) && ({row_reg, col_reg}<16'b0110101001100001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0110101001100001) && ({row_reg, col_reg}<16'b0110101001100011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110101001100011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110101001100100)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0110101001100101) && ({row_reg, col_reg}<16'b0110101001110001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0110101001110001) && ({row_reg, col_reg}<16'b0110101001110011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0110101001110011) && ({row_reg, col_reg}<16'b0110101001111010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110101001111010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0110101001111011) && ({row_reg, col_reg}<16'b0110101010001100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110101010001100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110101010001101) && ({row_reg, col_reg}<16'b0110101010001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110101010001111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110101010010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110101010010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110101010010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101010010011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110101010010100) && ({row_reg, col_reg}<16'b0110101010010111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110101010010111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110101010011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110101010011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101010011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110101010011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101010011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110101010011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110101010011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110101010011111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110101010100000) && ({row_reg, col_reg}<16'b0110101010100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101010100010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0110101010100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110101010100100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0110101010100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110101010100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0110101010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110101010101000) && ({row_reg, col_reg}<16'b0110101010101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110101010101010) && ({row_reg, col_reg}<16'b0110101010101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101010101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110101010101110) && ({row_reg, col_reg}<16'b0110101010110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110101010110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110101010110001) && ({row_reg, col_reg}<16'b0110101010110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110101010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110101010110101) && ({row_reg, col_reg}<16'b0110101010110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110101010110111) && ({row_reg, col_reg}<16'b0110101010111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110101010111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0110101010111100) && ({row_reg, col_reg}<16'b0110101010111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110101010111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110101011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101011000001) && ({row_reg, col_reg}<16'b0110101011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110101011000100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101011000101) && ({row_reg, col_reg}<16'b0110101011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101011010001) && ({row_reg, col_reg}<16'b0110101011110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110101011110111) && ({row_reg, col_reg}<16'b0110101011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110101011111001) && ({row_reg, col_reg}<16'b0110101011111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101011111011) && ({row_reg, col_reg}<16'b0110101011111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101011111110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}==16'b0110101011111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101100000000) && ({row_reg, col_reg}<16'b0110101100000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110101100000011) && ({row_reg, col_reg}<16'b0110101100000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101100000111) && ({row_reg, col_reg}<16'b0110101100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110101100001001) && ({row_reg, col_reg}<16'b0110101100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101100001101) && ({row_reg, col_reg}<16'b0110101100001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110101100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101100010000) && ({row_reg, col_reg}<16'b0110101100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101100010010) && ({row_reg, col_reg}<16'b0110101100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110101100100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101100100110) && ({row_reg, col_reg}<16'b0110101100101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110101100101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101100101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101100101110) && ({row_reg, col_reg}<16'b0110101100110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101100110001) && ({row_reg, col_reg}<16'b0110101100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110101100110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101100110100) && ({row_reg, col_reg}<16'b0110101100110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110101100110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110101100111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110101100111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110101100111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110101100111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110101100111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110101100111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110101100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101100111111) && ({row_reg, col_reg}<16'b0110101101000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110101101000010) && ({row_reg, col_reg}<16'b0110101101000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110101101000100) && ({row_reg, col_reg}<16'b0110101101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110101101000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110101101000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110101101001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110101101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110101101001100) && ({row_reg, col_reg}<16'b0110101101001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110101101001110) && ({row_reg, col_reg}<16'b0110101101010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101101010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110101101010100) && ({row_reg, col_reg}<16'b0110101101010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101101010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110101101010111) && ({row_reg, col_reg}<16'b0110101101011001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110101101011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110101101011010) && ({row_reg, col_reg}<16'b0110101101011100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110101101011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110101101011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110101101011110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110101101011111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110101101100000)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0110101101100001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110101101100010)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0110101101100011) && ({row_reg, col_reg}<16'b0110101101100101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110101101100101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0110101101100110) && ({row_reg, col_reg}<16'b0110101101110001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0110101101110001) && ({row_reg, col_reg}<16'b0110101101110011)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}>=16'b0110101101110011) && ({row_reg, col_reg}<16'b0110101101111001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110101101111001)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0110101101111010)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0110101101111011)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0110101101111100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0110101101111101) && ({row_reg, col_reg}<16'b0110101101111111)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=16'b0110101101111111) && ({row_reg, col_reg}<16'b0110101110001101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0110101110001101) && ({row_reg, col_reg}<16'b0110101110001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110101110001111) && ({row_reg, col_reg}<16'b0110101110010001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0110101110010001) && ({row_reg, col_reg}<16'b0110101110010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110101110010011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110101110010100) && ({row_reg, col_reg}<16'b0110101110010110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0110101110010110) && ({row_reg, col_reg}<16'b0110101110011000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110101110011000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110101110011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101110011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110101110011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101110011100) && ({row_reg, col_reg}<16'b0110101110011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110101110011110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110101110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101110100000) && ({row_reg, col_reg}<16'b0110101110100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110101110100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101110100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110101110100100) && ({row_reg, col_reg}<16'b0110101110100110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110101110100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110101110100111) && ({row_reg, col_reg}<16'b0110101110101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101110101010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0110101110101011) && ({row_reg, col_reg}<16'b0110101110101110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110101110101110) && ({row_reg, col_reg}<16'b0110101110110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110101110110000) && ({row_reg, col_reg}<16'b0110101110110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110101110110010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110101110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101110110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110101110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110101110110110) && ({row_reg, col_reg}<16'b0110101110111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110101110111000) && ({row_reg, col_reg}<16'b0110101110111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110101110111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110101110111101) && ({row_reg, col_reg}<16'b0110101111000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110101111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101111000001) && ({row_reg, col_reg}<16'b0110101111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110101111000100) && ({row_reg, col_reg}<16'b0110101111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101111000110) && ({row_reg, col_reg}<16'b0110101111001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101111001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101111001100) && ({row_reg, col_reg}<16'b0110101111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101111010001) && ({row_reg, col_reg}<16'b0110101111110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110101111110111) && ({row_reg, col_reg}<16'b0110101111111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110101111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110101111111010) && ({row_reg, col_reg}<16'b0110101111111100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0110101111111100) && ({row_reg, col_reg}<16'b0110110000000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110000000001) && ({row_reg, col_reg}<16'b0110110000000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110110000000011) && ({row_reg, col_reg}<16'b0110110000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110000000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110110000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110000000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110000001000) && ({row_reg, col_reg}<16'b0110110000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110000001101) && ({row_reg, col_reg}<16'b0110110000001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110000001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110000010000) && ({row_reg, col_reg}<16'b0110110000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110000010011) && ({row_reg, col_reg}<16'b0110110000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110000100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110000100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110110000100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110000101000) && ({row_reg, col_reg}<16'b0110110000101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110000101100) && ({row_reg, col_reg}<16'b0110110000101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110000101110) && ({row_reg, col_reg}<16'b0110110000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110000110001) && ({row_reg, col_reg}<16'b0110110000110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110000110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110110000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110110000110111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0110110000111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110110000111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110110000111010) && ({row_reg, col_reg}<16'b0110110000111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110000111100) && ({row_reg, col_reg}<16'b0110110000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110110000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110000111111) && ({row_reg, col_reg}<16'b0110110001000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110110001000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110110001000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110110001000110) && ({row_reg, col_reg}<16'b0110110001001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110110001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110110001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110110001001100) && ({row_reg, col_reg}<16'b0110110001001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110110001001110) && ({row_reg, col_reg}<16'b0110110001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110001010000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110110001010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110110001010010) && ({row_reg, col_reg}<16'b0110110001010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110110001010101) && ({row_reg, col_reg}<16'b0110110001010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110110001010111) && ({row_reg, col_reg}<16'b0110110001011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110110001011001) && ({row_reg, col_reg}<16'b0110110001011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110110001011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110110001011100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0110110001011101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0110110001011110)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0110110001011111) && ({row_reg, col_reg}<16'b0110110001100001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110110001100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110110001100010) && ({row_reg, col_reg}<16'b0110110001100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110110001100101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110110001100110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0110110001100111) && ({row_reg, col_reg}<16'b0110110001101111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110110001101111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110110001110000)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}>=16'b0110110001110001) && ({row_reg, col_reg}<16'b0110110001110011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0110110001110011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110110001110100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0110110001110101) && ({row_reg, col_reg}<16'b0110110001111000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110110001111000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110110001111001)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0110110001111010)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0110110001111011)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0110110001111100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0110110001111101) && ({row_reg, col_reg}<16'b0110110001111111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0110110001111111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110110010000000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0110110010000001) && ({row_reg, col_reg}<16'b0110110010010001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110110010010001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110110010010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110110010010011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110110010010100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0110110010010101) && ({row_reg, col_reg}<16'b0110110010010111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110110010010111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110110010011000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110110010011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110110010011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110010011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110010011100) && ({row_reg, col_reg}<16'b0110110010011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110010011110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110110010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110010100000) && ({row_reg, col_reg}<16'b0110110010100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110110010100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110110010100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110110010100100) && ({row_reg, col_reg}<16'b0110110010100110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110110010100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110110010100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110110010101000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110110010101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110110010101010) && ({row_reg, col_reg}<16'b0110110010101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110110010101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110010101101)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0110110010101110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110110010101111) && ({row_reg, col_reg}<16'b0110110010110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110110010110010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110110010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110010110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110110010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110010110110) && ({row_reg, col_reg}<16'b0110110010111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110110010111010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0110110010111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110110010111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110110010111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110010111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110110010111111) && ({row_reg, col_reg}<16'b0110110011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110011000001) && ({row_reg, col_reg}<16'b0110110011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110011000100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110110011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110110011000110) && ({row_reg, col_reg}<16'b0110110011001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110110011001100) && ({row_reg, col_reg}<16'b0110110011001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110011001111) && ({row_reg, col_reg}<16'b0110110011010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110011010001) && ({row_reg, col_reg}<16'b0110110011110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110110011110111) && ({row_reg, col_reg}<16'b0110110011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110110011111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110011111010) && ({row_reg, col_reg}<16'b0110110011111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110011111100) && ({row_reg, col_reg}<16'b0110110011111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110110011111110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}==16'b0110110011111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110110100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110100000001) && ({row_reg, col_reg}<16'b0110110100000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110110100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110100001000) && ({row_reg, col_reg}<16'b0110110100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110100001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110110100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110100010000) && ({row_reg, col_reg}<16'b0110110100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110100010011) && ({row_reg, col_reg}<16'b0110110100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110100100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110100100110) && ({row_reg, col_reg}<16'b0110110100101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110110100101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110100101100) && ({row_reg, col_reg}<16'b0110110100101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110100101110) && ({row_reg, col_reg}<16'b0110110100110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110100110001) && ({row_reg, col_reg}<16'b0110110100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110110100110100) && ({row_reg, col_reg}<16'b0110110100110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110110100110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110110100111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110110100111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110110100111010) && ({row_reg, col_reg}<16'b0110110100111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110110100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110100111111) && ({row_reg, col_reg}<16'b0110110101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110110101000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110110101000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110110101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110110101000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110101001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110110101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110110101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110110101001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110110101001101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0110110101001110) && ({row_reg, col_reg}<16'b0110110101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110101010000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110110101010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110110101010010) && ({row_reg, col_reg}<16'b0110110101010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110110101010101) && ({row_reg, col_reg}<16'b0110110101011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110110101011001) && ({row_reg, col_reg}<16'b0110110101011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110110101011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110101011100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0110110101011101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110110101011110)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0110110101011111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110110101100000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110110101100001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110110101100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110110101100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110110101100100) && ({row_reg, col_reg}<16'b0110110101100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110110101100110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110110101100111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110110101101000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110110101101001)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}>=16'b0110110101101010) && ({row_reg, col_reg}<16'b0110110101101100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110110101101100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110110101101101)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0110110101101110)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}>=16'b0110110101101111) && ({row_reg, col_reg}<16'b0110110101110001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110110101110001)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0110110101110010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0110110101110011)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0110110101110100)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}>=16'b0110110101110101) && ({row_reg, col_reg}<16'b0110110101110111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0110110101110111) && ({row_reg, col_reg}<16'b0110110101111001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110110101111001)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0110110101111010)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}>=16'b0110110101111011) && ({row_reg, col_reg}<16'b0110110101111101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110110101111101)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0110110101111110)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0110110101111111)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0110110110000000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0110110110000001) && ({row_reg, col_reg}<16'b0110110110000101)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0110110110000101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110110110000110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0110110110000111) && ({row_reg, col_reg}<16'b0110110110001010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110110110001010)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0110110110001011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110110110001100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0110110110001101) && ({row_reg, col_reg}<16'b0110110110010000)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0110110110010000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110110110010001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110110110010010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110110110010011) && ({row_reg, col_reg}<16'b0110110110010101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110110110010101) && ({row_reg, col_reg}<16'b0110110110010111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110110110010111) && ({row_reg, col_reg}<16'b0110110110011001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110110110011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110110110011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110110110011011) && ({row_reg, col_reg}<16'b0110110110011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110110011110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110110110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110110100000) && ({row_reg, col_reg}<16'b0110110110100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110110110100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110110100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110110110100100) && ({row_reg, col_reg}<16'b0110110110100110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110110110100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110110110100111) && ({row_reg, col_reg}<16'b0110110110101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110110110101010) && ({row_reg, col_reg}<16'b0110110110101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110110110101100) && ({row_reg, col_reg}<16'b0110110110101110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110110101110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0110110110101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110110110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110110110110001) && ({row_reg, col_reg}<16'b0110110110110011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110110110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110110110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110110110110101) && ({row_reg, col_reg}<16'b0110110110110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110110110111) && ({row_reg, col_reg}<16'b0110110110111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110110110111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110110110111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110110110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110110111110) && ({row_reg, col_reg}<16'b0110110111000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110111000001) && ({row_reg, col_reg}<16'b0110110111000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110110111000110) && ({row_reg, col_reg}<16'b0110110111001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110111001001) && ({row_reg, col_reg}<16'b0110110111001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110111001011) && ({row_reg, col_reg}<16'b0110110111001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110110111001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110110111001111) && ({row_reg, col_reg}<16'b0110110111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110111010001) && ({row_reg, col_reg}<16'b0110110111110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110111110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110111111000) && ({row_reg, col_reg}<16'b0110110111111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110110111111011)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0110110111111100) && ({row_reg, col_reg}<16'b0110111000000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111000000000) && ({row_reg, col_reg}<16'b0110111000000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111000000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110111000000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111000000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110111000000110) && ({row_reg, col_reg}<16'b0110111000001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111000001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110111000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111000001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110111000001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110111000001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110111000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111000010010) && ({row_reg, col_reg}<16'b0110111000100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110111000100110) && ({row_reg, col_reg}<16'b0110111000101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111000101000) && ({row_reg, col_reg}<16'b0110111000101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111000101100) && ({row_reg, col_reg}<16'b0110111000101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110111000101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111000101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110111000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111000110001) && ({row_reg, col_reg}<16'b0110111000110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110111000110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110111000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110111000110111) && ({row_reg, col_reg}<16'b0110111000111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111000111001) && ({row_reg, col_reg}<16'b0110111000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110111000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111000111111) && ({row_reg, col_reg}<16'b0110111001000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110111001000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110111001000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111001000110) && ({row_reg, col_reg}<16'b0110111001001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110111001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111001001010) && ({row_reg, col_reg}<16'b0110111001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110111001001100) && ({row_reg, col_reg}<16'b0110111001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111001001111) && ({row_reg, col_reg}<16'b0110111001010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110111001010011) && ({row_reg, col_reg}<16'b0110111001010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111001010111) && ({row_reg, col_reg}<16'b0110111001011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110111001011100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0110111001011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110111001011110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110111001011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111001100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110111001100001) && ({row_reg, col_reg}<16'b0110111001100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110111001100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110111001100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110111001100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0110111001100110) && ({row_reg, col_reg}<16'b0110111001101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110111001101000) && ({row_reg, col_reg}<16'b0110111001101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110111001101010) && ({row_reg, col_reg}<16'b0110111001101100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110111001101100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110111001101101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110111001101110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110111001101111) && ({row_reg, col_reg}<16'b0110111001110001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110111001110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111001110010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110111001110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110111001110100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110111001110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110111001110110) && ({row_reg, col_reg}<16'b0110111001111010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110111001111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110111001111011) && ({row_reg, col_reg}<16'b0110111001111101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110111001111101) && ({row_reg, col_reg}<16'b0110111010000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110111010000000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0110111010000001) && ({row_reg, col_reg}<16'b0110111010000011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110111010000011) && ({row_reg, col_reg}<16'b0110111010000101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0110111010000101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110111010000110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110111010000111) && ({row_reg, col_reg}<16'b0110111010001010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110111010001010) && ({row_reg, col_reg}<16'b0110111010001100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110111010001100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110111010001101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0110111010001110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0110111010001111) && ({row_reg, col_reg}<16'b0110111010010001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110111010010001) && ({row_reg, col_reg}<16'b0110111010010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111010010111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110111010011000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110111010011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111010011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110111010011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111010011100) && ({row_reg, col_reg}<16'b0110111010011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110111010011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111010011111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110111010100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110111010100001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0110111010100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110111010100011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110111010100100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110111010100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110111010100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0110111010100111) && ({row_reg, col_reg}<16'b0110111010101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110111010101001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110111010101010) && ({row_reg, col_reg}<16'b0110111010101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110111010101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110111010101101) && ({row_reg, col_reg}<16'b0110111010110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111010110000) && ({row_reg, col_reg}<16'b0110111010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110111010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110111010110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110111010110101) && ({row_reg, col_reg}<16'b0110111010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111010111000) && ({row_reg, col_reg}<16'b0110111010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111010111010) && ({row_reg, col_reg}<16'b0110111011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111011000001) && ({row_reg, col_reg}<16'b0110111011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110111011000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111011000110) && ({row_reg, col_reg}<16'b0110111011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110111011001010)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==16'b0110111011001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111011001100) && ({row_reg, col_reg}<16'b0110111011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111011001111) && ({row_reg, col_reg}<16'b0110111011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111011010001) && ({row_reg, col_reg}<16'b0110111011110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110111011110100) && ({row_reg, col_reg}<16'b0110111011110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111011110110) && ({row_reg, col_reg}<16'b0110111011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110111011111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111011111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111011111101) && ({row_reg, col_reg}<16'b0110111011111111)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}==16'b0110111011111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111100000000) && ({row_reg, col_reg}<16'b0110111100001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111100001011) && ({row_reg, col_reg}<16'b0110111100001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111100001101) && ({row_reg, col_reg}<16'b0110111100001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110111100001111) && ({row_reg, col_reg}<16'b0110111100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111100010010) && ({row_reg, col_reg}<16'b0110111100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110111100100110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111100100111) && ({row_reg, col_reg}<16'b0110111100101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111100101010) && ({row_reg, col_reg}<16'b0110111100101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110111100101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111100101110) && ({row_reg, col_reg}<16'b0110111100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110111100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111100110001) && ({row_reg, col_reg}<16'b0110111100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110111100110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110111100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111100110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110111100110111) && ({row_reg, col_reg}<16'b0110111100111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110111100111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110111100111010) && ({row_reg, col_reg}<16'b0110111100111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111100111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110111100111101) && ({row_reg, col_reg}<16'b0110111100111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111100111111) && ({row_reg, col_reg}<16'b0110111101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110111101000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110111101000101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0110111101000110) && ({row_reg, col_reg}<16'b0110111101001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110111101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110111101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111101001100) && ({row_reg, col_reg}<16'b0110111101001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110111101001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111101001111) && ({row_reg, col_reg}<16'b0110111101010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110111101010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110111101010100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0110111101010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110111101010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111101010111) && ({row_reg, col_reg}<16'b0110111101011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110111101011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111101011010) && ({row_reg, col_reg}<16'b0110111101011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110111101011100) && ({row_reg, col_reg}<16'b0110111101011110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110111101011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111101011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110111101100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110111101100001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110111101100010) && ({row_reg, col_reg}<16'b0110111101100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111101100110) && ({row_reg, col_reg}<16'b0110111101101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110111101101000) && ({row_reg, col_reg}<16'b0110111101101010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110111101101010) && ({row_reg, col_reg}<16'b0110111101101100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0110111101101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111101101101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110111101101110) && ({row_reg, col_reg}<16'b0110111101110001)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0110111101110001) && ({row_reg, col_reg}<16'b0110111101110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110111101110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111101110100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110111101110101) && ({row_reg, col_reg}<16'b0110111101111010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0110111101111010) && ({row_reg, col_reg}<16'b0110111101111100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110111101111100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0110111101111101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110111101111110) && ({row_reg, col_reg}<16'b0110111110000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111110000101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110111110000110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0110111110000111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110111110001000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111110001001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110111110001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110111110001011) && ({row_reg, col_reg}<16'b0110111110001101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110111110001101) && ({row_reg, col_reg}<16'b0110111110010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111110010000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110111110010001) && ({row_reg, col_reg}<16'b0110111110010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111110010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110111110010100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110111110010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111110010110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110111110010111) && ({row_reg, col_reg}<16'b0110111110011001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0110111110011001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110111110011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110111110011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110111110011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111110011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110111110011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111110011111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110111110100000) && ({row_reg, col_reg}<16'b0110111110100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110111110100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110111110100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111110100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110111110100101) && ({row_reg, col_reg}<16'b0110111110100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110111110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111110101001) && ({row_reg, col_reg}<16'b0110111110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111110101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110111110101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111110101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111110101110) && ({row_reg, col_reg}<16'b0110111110110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111110110001) && ({row_reg, col_reg}<16'b0110111110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110111110110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110111110110100) && ({row_reg, col_reg}<16'b0110111110110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111110110110) && ({row_reg, col_reg}<16'b0110111110111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111110111001) && ({row_reg, col_reg}<16'b0110111110111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110111110111011) && ({row_reg, col_reg}<16'b0110111110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110111110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111110111110) && ({row_reg, col_reg}<16'b0110111111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110111111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111111000001) && ({row_reg, col_reg}<16'b0110111111000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110111111000101) && ({row_reg, col_reg}<16'b0110111111000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111111000111) && ({row_reg, col_reg}<16'b0110111111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111111001001) && ({row_reg, col_reg}<16'b0110111111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111111001011) && ({row_reg, col_reg}<16'b0110111111001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111111001111) && ({row_reg, col_reg}<16'b0110111111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111111010001) && ({row_reg, col_reg}<16'b0110111111110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110111111110100) && ({row_reg, col_reg}<16'b0110111111110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111111110110) && ({row_reg, col_reg}<16'b0110111111111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111111111010) && ({row_reg, col_reg}<16'b0110111111111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111111111100) && ({row_reg, col_reg}<16'b0110111111111111)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}==16'b0110111111111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000000000000) && ({row_reg, col_reg}<16'b0111000000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000000001100) && ({row_reg, col_reg}<16'b0111000000001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000000001110) && ({row_reg, col_reg}<16'b0111000000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000000010010) && ({row_reg, col_reg}<16'b0111000000100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000000100110) && ({row_reg, col_reg}<16'b0111000000101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111000000101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000000101001) && ({row_reg, col_reg}<16'b0111000000101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000000101011) && ({row_reg, col_reg}<16'b0111000000101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000000101101) && ({row_reg, col_reg}<16'b0111000000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000000110001) && ({row_reg, col_reg}<16'b0111000000110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111000000110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111000000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000000110110) && ({row_reg, col_reg}<16'b0111000000111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000000111001) && ({row_reg, col_reg}<16'b0111000000111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000000111100) && ({row_reg, col_reg}<16'b0111000000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111000000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000000111111) && ({row_reg, col_reg}<16'b0111000001000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000001000100) && ({row_reg, col_reg}<16'b0111000001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111000001000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111000001000111) && ({row_reg, col_reg}<16'b0111000001001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111000001001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111000001001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000001001011) && ({row_reg, col_reg}<16'b0111000001001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111000001001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000001001110) && ({row_reg, col_reg}<16'b0111000001010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111000001010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111000001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111000001010101)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0111000001010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0111000001010111) && ({row_reg, col_reg}<16'b0111000001011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111000001011011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111000001011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111000001011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111000001011110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0111000001011111) && ({row_reg, col_reg}<16'b0111000001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111000001100010) && ({row_reg, col_reg}<16'b0111000001100100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0111000001100100) && ({row_reg, col_reg}<16'b0111000010010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111000010010001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111000010010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111000010010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111000010010100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111000010010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111000010010110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0111000010010111) && ({row_reg, col_reg}<16'b0111000010011001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0111000010011001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111000010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111000010011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111000010011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111000010011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111000010011110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111000010011111) && ({row_reg, col_reg}<16'b0111000010100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111000010100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111000010100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0111000010100100) && ({row_reg, col_reg}<16'b0111000010100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111000010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111000010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111000010101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000010101010) && ({row_reg, col_reg}<16'b0111000010101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111000010101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000010101110) && ({row_reg, col_reg}<16'b0111000010110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000010110000) && ({row_reg, col_reg}<16'b0111000010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111000010110011) && ({row_reg, col_reg}<16'b0111000010110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111000010110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000010110110) && ({row_reg, col_reg}<16'b0111000010111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000010111001) && ({row_reg, col_reg}<16'b0111000010111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111000010111011) && ({row_reg, col_reg}<16'b0111000010111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111000010111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111000010111111) && ({row_reg, col_reg}<16'b0111000011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000011000001) && ({row_reg, col_reg}<16'b0111000011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000011000101) && ({row_reg, col_reg}<16'b0111000011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111000011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111000011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111000011001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111000011001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111000011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000011001111) && ({row_reg, col_reg}<16'b0111000011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000011010001) && ({row_reg, col_reg}<16'b0111000011110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000011110100) && ({row_reg, col_reg}<16'b0111000011110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000011110110) && ({row_reg, col_reg}<16'b0111000011111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111000011111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111000011111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0111000011111100) && ({row_reg, col_reg}<16'b0111000100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000100000000) && ({row_reg, col_reg}<16'b0111000100000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111000100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000100001000) && ({row_reg, col_reg}<16'b0111000100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000100001101) && ({row_reg, col_reg}<16'b0111000100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000100001111) && ({row_reg, col_reg}<16'b0111000100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000100010010) && ({row_reg, col_reg}<16'b0111000100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111000100100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000100100110) && ({row_reg, col_reg}<16'b0111000100101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111000100101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000100101011) && ({row_reg, col_reg}<16'b0111000100101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000100101101) && ({row_reg, col_reg}<16'b0111000100110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000100110001) && ({row_reg, col_reg}<16'b0111000100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111000100110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111000100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000100110110) && ({row_reg, col_reg}<16'b0111000100111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000100111001) && ({row_reg, col_reg}<16'b0111000100111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000100111100) && ({row_reg, col_reg}<16'b0111000100111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111000100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000100111111) && ({row_reg, col_reg}<16'b0111000101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111000101000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111000101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111000101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111000101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111000101000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111000101001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111000101001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111000101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111000101001011) && ({row_reg, col_reg}<16'b0111000101001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111000101001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000101001110) && ({row_reg, col_reg}<16'b0111000101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111000101010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111000101010001) && ({row_reg, col_reg}<16'b0111000101010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111000101010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111000101010100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0111000101010101)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0111000101010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0111000101010111) && ({row_reg, col_reg}<16'b0111000101011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111000101011100) && ({row_reg, col_reg}<16'b0111000110010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111000110010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111000110010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111000110010101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111000110010110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0111000110010111) && ({row_reg, col_reg}<16'b0111000110011001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0111000110011001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111000110011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0111000110011011) && ({row_reg, col_reg}<16'b0111000110011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111000110011110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111000110011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000110100000) && ({row_reg, col_reg}<16'b0111000110100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111000110100011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0111000110100100) && ({row_reg, col_reg}<16'b0111000110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111000110100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0111000110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111000110101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000110101001) && ({row_reg, col_reg}<16'b0111000110101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111000110101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111000110101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111000110101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000110110000) && ({row_reg, col_reg}<16'b0111000110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111000110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111000110110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111000110110101) && ({row_reg, col_reg}<16'b0111000110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000110111000) && ({row_reg, col_reg}<16'b0111000110111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111000110111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111000110111011) && ({row_reg, col_reg}<16'b0111000110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000110111101) && ({row_reg, col_reg}<16'b0111000110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111000110111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111000111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000111000001) && ({row_reg, col_reg}<16'b0111000111000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111000111000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000111000110) && ({row_reg, col_reg}<16'b0111000111001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111000111001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000111001100) && ({row_reg, col_reg}<16'b0111000111001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000111001111) && ({row_reg, col_reg}<16'b0111000111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000111010001) && ({row_reg, col_reg}<16'b0111000111110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000111110100) && ({row_reg, col_reg}<16'b0111000111110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000111110111) && ({row_reg, col_reg}<16'b0111000111111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111000111111010)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0111000111111011) && ({row_reg, col_reg}<16'b0111001000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111001000000000) && ({row_reg, col_reg}<16'b0111001000000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001000000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001000001000) && ({row_reg, col_reg}<16'b0111001000001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001000001010) && ({row_reg, col_reg}<16'b0111001000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111001000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001000001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111001000001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001000001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001000010000) && ({row_reg, col_reg}<16'b0111001000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001000010011) && ({row_reg, col_reg}<16'b0111001000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001000100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001000100110) && ({row_reg, col_reg}<16'b0111001000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001000110001) && ({row_reg, col_reg}<16'b0111001000110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001000110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111001000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001000110110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0111001000110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001000111001) && ({row_reg, col_reg}<16'b0111001000111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001000111100) && ({row_reg, col_reg}<16'b0111001000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111001000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001000111111) && ({row_reg, col_reg}<16'b0111001001000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111001001000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111001001000100) && ({row_reg, col_reg}<16'b0111001001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001001000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111001001000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001001001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111001001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111001001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111001001001100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111001001001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111001001001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111001001001111) && ({row_reg, col_reg}<16'b0111001001010001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111001001010001) && ({row_reg, col_reg}<16'b0111001001010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111001001010101) && ({row_reg, col_reg}<16'b0111001001010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0111001001010111) && ({row_reg, col_reg}<16'b0111001001011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001001011001)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0111001001011010) && ({row_reg, col_reg}<16'b0111001001011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001001011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001001011101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111001001011110) && ({row_reg, col_reg}<16'b0111001001100000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111001001100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001001100001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111001001100010) && ({row_reg, col_reg}<16'b0111001001100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111001001100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111001001100110) && ({row_reg, col_reg}<16'b0111001001101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001001101001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111001001101010) && ({row_reg, col_reg}<16'b0111001001101100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111001001101100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111001001101101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111001001101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001001101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111001001110000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111001001110001) && ({row_reg, col_reg}<16'b0111001001111001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111001001111001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111001001111010) && ({row_reg, col_reg}<16'b0111001001111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111001001111100) && ({row_reg, col_reg}<16'b0111001001111111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111001001111111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111001010000000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111001010000001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111001010000010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111001010000011) && ({row_reg, col_reg}<16'b0111001010001010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111001010001010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111001010001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001010001100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111001010001101) && ({row_reg, col_reg}<16'b0111001010001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111001010001111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111001010010000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111001010010001) && ({row_reg, col_reg}<16'b0111001010010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001010010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111001010010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001010010101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111001010010110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0111001010010111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0111001010011000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0111001010011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001010011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001010011011) && ({row_reg, col_reg}<16'b0111001010011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001010011110) && ({row_reg, col_reg}<16'b0111001010100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001010100000) && ({row_reg, col_reg}<16'b0111001010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001010100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0111001010100100) && ({row_reg, col_reg}<16'b0111001010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111001010100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0111001010100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111001010101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001010101001) && ({row_reg, col_reg}<16'b0111001010101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001010101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111001010101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001010101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111001010110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001010110001) && ({row_reg, col_reg}<16'b0111001010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111001010110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111001010110101) && ({row_reg, col_reg}<16'b0111001010110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111001010110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111001010111000) && ({row_reg, col_reg}<16'b0111001010111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0111001010111010) && ({row_reg, col_reg}<16'b0111001010111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111001010111100) && ({row_reg, col_reg}<16'b0111001010111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111001010111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111001011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001011000001) && ({row_reg, col_reg}<16'b0111001011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001011000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001011000110) && ({row_reg, col_reg}<16'b0111001011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001011001010) && ({row_reg, col_reg}<16'b0111001011001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001011001100) && ({row_reg, col_reg}<16'b0111001011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001011010001) && ({row_reg, col_reg}<16'b0111001011110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001011110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001011110101) && ({row_reg, col_reg}<16'b0111001011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111001011111000) && ({row_reg, col_reg}<16'b0111001011111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001011111010)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0111001011111011) && ({row_reg, col_reg}<16'b0111001100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111001100000000) && ({row_reg, col_reg}<16'b0111001100001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001100001010) && ({row_reg, col_reg}<16'b0111001100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111001100001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001100001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111001100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001100010000) && ({row_reg, col_reg}<16'b0111001100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001100010011) && ({row_reg, col_reg}<16'b0111001100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111001100100100) && ({row_reg, col_reg}<16'b0111001100100110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001100100110) && ({row_reg, col_reg}<16'b0111001100101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001100101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001100101111) && ({row_reg, col_reg}<16'b0111001100110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001100110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001100110010) && ({row_reg, col_reg}<16'b0111001100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111001100110100) && ({row_reg, col_reg}<16'b0111001100110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001100110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111001100110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001100111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001100111001) && ({row_reg, col_reg}<16'b0111001100111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001100111100) && ({row_reg, col_reg}<16'b0111001100111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111001100111111) && ({row_reg, col_reg}<16'b0111001101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111001101000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111001101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111001101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001101000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111001101000111) && ({row_reg, col_reg}<16'b0111001101001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111001101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001101001010) && ({row_reg, col_reg}<16'b0111001101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111001101001100) && ({row_reg, col_reg}<16'b0111001101001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001101001110) && ({row_reg, col_reg}<16'b0111001101011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111001101011001) && ({row_reg, col_reg}<16'b0111001101011011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111001101011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001101011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001101011101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111001101011110) && ({row_reg, col_reg}<16'b0111001101100000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111001101100000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111001101100001) && ({row_reg, col_reg}<16'b0111001101100110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0111001101100110) && ({row_reg, col_reg}<16'b0111001101101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001101101001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111001101101010) && ({row_reg, col_reg}<16'b0111001101101100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111001101101100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111001101101101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111001101101110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111001101101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111001101110000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111001101110001) && ({row_reg, col_reg}<16'b0111001101111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111001101111010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111001101111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111001101111100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111001101111101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111001101111110) && ({row_reg, col_reg}<16'b0111001110000001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111001110000001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111001110000010) && ({row_reg, col_reg}<16'b0111001110001011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111001110001011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111001110001100) && ({row_reg, col_reg}<16'b0111001110001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0111001110001111) && ({row_reg, col_reg}<16'b0111001110010001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111001110010001) && ({row_reg, col_reg}<16'b0111001110010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001110010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111001110010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001110010101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111001110010110) && ({row_reg, col_reg}<16'b0111001110011000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0111001110011000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111001110011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001110011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111001110011011) && ({row_reg, col_reg}<16'b0111001110011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111001110011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111001110011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001110100000) && ({row_reg, col_reg}<16'b0111001110100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001110100011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0111001110100100) && ({row_reg, col_reg}<16'b0111001110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111001110100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0111001110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111001110101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111001110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001110101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001110101011) && ({row_reg, col_reg}<16'b0111001110101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001110101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111001110101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001110110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111001110110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111001110110010) && ({row_reg, col_reg}<16'b0111001110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001110110100) && ({row_reg, col_reg}<16'b0111001110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001110111000) && ({row_reg, col_reg}<16'b0111001110111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111001110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111001110111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111001110111100) && ({row_reg, col_reg}<16'b0111001110111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111001110111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111001111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001111000001) && ({row_reg, col_reg}<16'b0111001111000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001111000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001111000110) && ({row_reg, col_reg}<16'b0111001111001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001111001010) && ({row_reg, col_reg}<16'b0111001111001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001111001100) && ({row_reg, col_reg}<16'b0111001111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001111001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001111001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001111010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001111010001) && ({row_reg, col_reg}<16'b0111001111110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001111110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001111110101) && ({row_reg, col_reg}<16'b0111001111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001111111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111001111111010)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0111001111111011) && ({row_reg, col_reg}<16'b0111010000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111010000000000) && ({row_reg, col_reg}<16'b0111010000001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010000001001) && ({row_reg, col_reg}<16'b0111010000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111010000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010000001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111010000001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111010000001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010000010000) && ({row_reg, col_reg}<16'b0111010000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010000010010) && ({row_reg, col_reg}<16'b0111010000100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111010000100100) && ({row_reg, col_reg}<16'b0111010000100110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010000100110) && ({row_reg, col_reg}<16'b0111010000101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010000101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111010000101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010000110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010000110001) && ({row_reg, col_reg}<16'b0111010000110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111010000110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010000110100) && ({row_reg, col_reg}<16'b0111010000110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111010000110111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0111010000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111010000111001) && ({row_reg, col_reg}<16'b0111010000111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111010000111100) && ({row_reg, col_reg}<16'b0111010000111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111010000111111) && ({row_reg, col_reg}<16'b0111010001000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111010001000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111010001000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111010001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111010001000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111010001000111) && ({row_reg, col_reg}<16'b0111010001001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111010001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111010001001010) && ({row_reg, col_reg}<16'b0111010001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111010001001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111010001001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111010001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111010001001111) && ({row_reg, col_reg}<16'b0111010001010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111010001010010) && ({row_reg, col_reg}<16'b0111010001010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111010001010101) && ({row_reg, col_reg}<16'b0111010001011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111010001011001)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0111010001011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111010001011011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111010001011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111010001011101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111010001011110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111010001011111) && ({row_reg, col_reg}<16'b0111010001100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111010001100100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111010001100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111010001100110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111010001100111) && ({row_reg, col_reg}<16'b0111010001101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111010001101110) && ({row_reg, col_reg}<16'b0111010001110001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111010001110001) && ({row_reg, col_reg}<16'b0111010001111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111010001111010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111010001111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111010001111100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111010001111101) && ({row_reg, col_reg}<16'b0111010010000001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0111010010000001) && ({row_reg, col_reg}<16'b0111010010000011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111010010000011) && ({row_reg, col_reg}<16'b0111010010000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0111010010000110) && ({row_reg, col_reg}<16'b0111010010001010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111010010001010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111010010001011) && ({row_reg, col_reg}<16'b0111010010001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111010010001101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111010010001110) && ({row_reg, col_reg}<16'b0111010010010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111010010010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111010010010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111010010010101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0111010010010110) && ({row_reg, col_reg}<16'b0111010010011000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0111010010011000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0111010010011001) && ({row_reg, col_reg}<16'b0111010010011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111010010011011) && ({row_reg, col_reg}<16'b0111010010011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111010010011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111010010100000) && ({row_reg, col_reg}<16'b0111010010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111010010100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0111010010100100) && ({row_reg, col_reg}<16'b0111010010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111010010100110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111010010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111010010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111010010101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111010010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010010101011) && ({row_reg, col_reg}<16'b0111010010101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111010010101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111010010101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010010101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111010010110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111010010110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111010010110010)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}==16'b0111010010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111010010110100) && ({row_reg, col_reg}<16'b0111010010110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111010010110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111010010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111010010111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111010010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111010010111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111010010111100) && ({row_reg, col_reg}<16'b0111010010111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111010010111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111010011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010011000001) && ({row_reg, col_reg}<16'b0111010011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111010011000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010011000110) && ({row_reg, col_reg}<16'b0111010011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010011001001) && ({row_reg, col_reg}<16'b0111010011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111010011001011) && ({row_reg, col_reg}<16'b0111010011001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010011001101) && ({row_reg, col_reg}<16'b0111010011001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111010011001111) && ({row_reg, col_reg}<16'b0111010011010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010011010001) && ({row_reg, col_reg}<16'b0111010011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111010011111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111010011111010)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0111010011111011) && ({row_reg, col_reg}<16'b0111010100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111010100000000) && ({row_reg, col_reg}<16'b0111010100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111010100000010) && ({row_reg, col_reg}<16'b0111010100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010100000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010100000111) && ({row_reg, col_reg}<16'b0111010100001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010100001001) && ({row_reg, col_reg}<16'b0111010100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111010100001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010100001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111010100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111010100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111010100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010100010010) && ({row_reg, col_reg}<16'b0111010100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111010100100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010100100110) && ({row_reg, col_reg}<16'b0111010100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010100110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111010100110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111010100110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010100110011) && ({row_reg, col_reg}<16'b0111010100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010100110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111010100110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111010100110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111010100111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111010100111001) && ({row_reg, col_reg}<16'b0111010100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111010100111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010100111100) && ({row_reg, col_reg}<16'b0111010100111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111010100111111) && ({row_reg, col_reg}<16'b0111010101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111010101000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111010101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111010101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111010101000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111010101000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111010101001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111010101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111010101001010) && ({row_reg, col_reg}<16'b0111010101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111010101001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111010101001101) && ({row_reg, col_reg}<16'b0111010101001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111010101001111) && ({row_reg, col_reg}<16'b0111010101010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111010101010011) && ({row_reg, col_reg}<16'b0111010101010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0111010101010101) && ({row_reg, col_reg}<16'b0111010101011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111010101011001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0111010101011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0111010101011011) && ({row_reg, col_reg}<16'b0111010101011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111010101011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111010101011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111010101100000) && ({row_reg, col_reg}<16'b0111010101100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0111010101100100) && ({row_reg, col_reg}<16'b0111010101100111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111010101100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111010101101000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111010101101001) && ({row_reg, col_reg}<16'b0111010101101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111010101101011) && ({row_reg, col_reg}<16'b0111010101101101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111010101101101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111010101101110) && ({row_reg, col_reg}<16'b0111010101110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111010101110110) && ({row_reg, col_reg}<16'b0111010101111000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111010101111000) && ({row_reg, col_reg}<16'b0111010101111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111010101111010) && ({row_reg, col_reg}<16'b0111010101111100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111010101111100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111010101111101) && ({row_reg, col_reg}<16'b0111010110000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111010110000000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111010110000001) && ({row_reg, col_reg}<16'b0111010110000011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111010110000011) && ({row_reg, col_reg}<16'b0111010110001010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111010110001010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111010110001011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111010110001100) && ({row_reg, col_reg}<16'b0111010110001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111010110001110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111010110001111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111010110010000) && ({row_reg, col_reg}<16'b0111010110010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111010110010100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0111010110010101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0111010110010110)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0111010110010111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0111010110011000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0111010110011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111010110011010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0111010110011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111010110011100) && ({row_reg, col_reg}<16'b0111010110011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111010110011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111010110100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111010110100001) && ({row_reg, col_reg}<16'b0111010110100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111010110100011) && ({row_reg, col_reg}<16'b0111010110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111010110100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111010110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111010110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111010110101001) && ({row_reg, col_reg}<16'b0111010110101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111010110101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010110101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111010110101110) && ({row_reg, col_reg}<16'b0111010110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111010110110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111010110110101) && ({row_reg, col_reg}<16'b0111010110110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111010110110111) && ({row_reg, col_reg}<16'b0111010110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111010110111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111010111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010111000001) && ({row_reg, col_reg}<16'b0111010111000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111010111000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010111000110) && ({row_reg, col_reg}<16'b0111010111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010111001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111010111001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010111001011) && ({row_reg, col_reg}<16'b0111010111001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010111001101) && ({row_reg, col_reg}<16'b0111010111001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111010111001111) && ({row_reg, col_reg}<16'b0111010111010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010111010001) && ({row_reg, col_reg}<16'b0111010111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111010111111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111010111111010)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0111010111111011) && ({row_reg, col_reg}<16'b0111011000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111011000000000) && ({row_reg, col_reg}<16'b0111011000000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011000000010) && ({row_reg, col_reg}<16'b0111011000001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011000001010) && ({row_reg, col_reg}<16'b0111011000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011000001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111011000001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111011000001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111011000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011000010010) && ({row_reg, col_reg}<16'b0111011000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111011000100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011000100110) && ({row_reg, col_reg}<16'b0111011000101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011000101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111011000101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011000101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011000101100) && ({row_reg, col_reg}<16'b0111011000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011000110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111011000110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111011000110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111011000110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011000110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111011000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111011000110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111011000111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111011000111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011000111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011000111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111011000111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111011000111101) && ({row_reg, col_reg}<16'b0111011000111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111011000111111) && ({row_reg, col_reg}<16'b0111011001000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011001000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111011001000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111011001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111011001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111011001000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011001001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111011001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111011001001010) && ({row_reg, col_reg}<16'b0111011001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111011001001100) && ({row_reg, col_reg}<16'b0111011001010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111011001010000) && ({row_reg, col_reg}<16'b0111011001010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111011001010010) && ({row_reg, col_reg}<16'b0111011001010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111011001010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0111011001010110) && ({row_reg, col_reg}<16'b0111011001011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111011001011001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0111011001011010) && ({row_reg, col_reg}<16'b0111011001011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111011001011100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111011001011101) && ({row_reg, col_reg}<16'b0111011001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111011001011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111011001100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111011001100001) && ({row_reg, col_reg}<16'b0111011001100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111011001100100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111011001100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111011001100110) && ({row_reg, col_reg}<16'b0111011001101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111011001101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111011001101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111011001101010) && ({row_reg, col_reg}<16'b0111011001110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111011001110001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111011001110010) && ({row_reg, col_reg}<16'b0111011001111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111011001111101) && ({row_reg, col_reg}<16'b0111011001111111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111011001111111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111011010000000) && ({row_reg, col_reg}<16'b0111011010000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111011010000101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111011010000110) && ({row_reg, col_reg}<16'b0111011010001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111011010001100) && ({row_reg, col_reg}<16'b0111011010001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111011010001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111011010001111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111011010010000) && ({row_reg, col_reg}<16'b0111011010010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111011010010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111011010010011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0111011010010100)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0111011010010101) && ({row_reg, col_reg}<16'b0111011010011000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0111011010011000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0111011010011001) && ({row_reg, col_reg}<16'b0111011010011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111011010011011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111011010011100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=16'b0111011010011101) && ({row_reg, col_reg}<16'b0111011010100000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0111011010100000) && ({row_reg, col_reg}<16'b0111011010100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111011010100011) && ({row_reg, col_reg}<16'b0111011010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111011010100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111011010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111011010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111011010101001) && ({row_reg, col_reg}<16'b0111011010101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011010101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111011010101110) && ({row_reg, col_reg}<16'b0111011010110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111011010110001) && ({row_reg, col_reg}<16'b0111011010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111011010110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111011010110101) && ({row_reg, col_reg}<16'b0111011010110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011010110111) && ({row_reg, col_reg}<16'b0111011010111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111011010111001) && ({row_reg, col_reg}<16'b0111011010111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011010111011) && ({row_reg, col_reg}<16'b0111011010111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111011010111101) && ({row_reg, col_reg}<16'b0111011011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011011000001) && ({row_reg, col_reg}<16'b0111011011000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111011011000110) && ({row_reg, col_reg}<16'b0111011011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011011001010) && ({row_reg, col_reg}<16'b0111011011010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011011010001) && ({row_reg, col_reg}<16'b0111011011110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111011011110001) && ({row_reg, col_reg}<16'b0111011011110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011011110110) && ({row_reg, col_reg}<16'b0111011011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111011011111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111011011111010)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0111011011111011) && ({row_reg, col_reg}<16'b0111011100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111011100000000) && ({row_reg, col_reg}<16'b0111011100000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011100000011) && ({row_reg, col_reg}<16'b0111011100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011100001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111011100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111011100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111011100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011100010010) && ({row_reg, col_reg}<16'b0111011100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111011100100110) && ({row_reg, col_reg}<16'b0111011100101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011100101001) && ({row_reg, col_reg}<16'b0111011100101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011100101011) && ({row_reg, col_reg}<16'b0111011100110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011100110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111011100110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111011100110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011100110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111011100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011100110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111011100111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111011100111001) && ({row_reg, col_reg}<16'b0111011100111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111011100111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111011100111101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0111011100111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111011100111111) && ({row_reg, col_reg}<16'b0111011101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011101000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111011101000100) && ({row_reg, col_reg}<16'b0111011101000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111011101000111) && ({row_reg, col_reg}<16'b0111011101001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111011101001001) && ({row_reg, col_reg}<16'b0111011101001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111011101001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111011101001101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0111011101001110) && ({row_reg, col_reg}<16'b0111011101010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111011101010000) && ({row_reg, col_reg}<16'b0111011101010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111011101010010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111011101010011) && ({row_reg, col_reg}<16'b0111011101010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111011101010101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0111011101010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111011101010111) && ({row_reg, col_reg}<16'b0111011101011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111011101011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111011101011010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111011101011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111011101011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111011101011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111011101011110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111011101011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111011101100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111011101100001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111011101100010) && ({row_reg, col_reg}<16'b0111011101101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111011101101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111011101101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111011101101010) && ({row_reg, col_reg}<16'b0111011101101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111011101101100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111011101101101) && ({row_reg, col_reg}<16'b0111011101110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111011101110011) && ({row_reg, col_reg}<16'b0111011101110101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111011101110101) && ({row_reg, col_reg}<16'b0111011101110111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111011101110111) && ({row_reg, col_reg}<16'b0111011101111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111011101111010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111011101111011) && ({row_reg, col_reg}<16'b0111011101111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111011101111111) && ({row_reg, col_reg}<16'b0111011110000001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111011110000001) && ({row_reg, col_reg}<16'b0111011110000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111011110000011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111011110000100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111011110000101) && ({row_reg, col_reg}<16'b0111011110001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111011110001010) && ({row_reg, col_reg}<16'b0111011110001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111011110001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111011110001101) && ({row_reg, col_reg}<16'b0111011110001111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111011110001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111011110010000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111011110010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111011110010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111011110010011)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0111011110010100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111011110010101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0111011110010110)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0111011110010111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0111011110011000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0111011110011001) && ({row_reg, col_reg}<16'b0111011110011101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111011110011101) && ({row_reg, col_reg}<16'b0111011110100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111011110100011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0111011110100100) && ({row_reg, col_reg}<16'b0111011110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111011110100110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0111011110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111011110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111011110101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011110101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111011110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011110101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011110101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111011110101110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111011110101111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111011110110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111011110110001) && ({row_reg, col_reg}<16'b0111011110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111011110110011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0111011110110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111011110110101) && ({row_reg, col_reg}<16'b0111011110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011110111110) && ({row_reg, col_reg}<16'b0111011111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011111000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011111000010) && ({row_reg, col_reg}<16'b0111011111000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111011111000110) && ({row_reg, col_reg}<16'b0111011111001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011111001010) && ({row_reg, col_reg}<16'b0111011111001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011111001100) && ({row_reg, col_reg}<16'b0111011111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011111001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111011111001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011111010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011111010001) && ({row_reg, col_reg}<16'b0111011111110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111011111110000) && ({row_reg, col_reg}<16'b0111011111110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011111110011) && ({row_reg, col_reg}<16'b0111011111110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011111110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011111110111) && ({row_reg, col_reg}<16'b0111011111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111011111111001) && ({row_reg, col_reg}<16'b0111011111111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011111111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0111011111111100) && ({row_reg, col_reg}<16'b0111100000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111100000000000) && ({row_reg, col_reg}<16'b0111100000000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100000000011) && ({row_reg, col_reg}<16'b0111100000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100000000110) && ({row_reg, col_reg}<16'b0111100000001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111100000001000) && ({row_reg, col_reg}<16'b0111100000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111100000001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111100000001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111100000001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111100000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111100000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111100000010010) && ({row_reg, col_reg}<16'b0111100000100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111100000100110) && ({row_reg, col_reg}<16'b0111100000101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100000101010) && ({row_reg, col_reg}<16'b0111100000101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100000101100) && ({row_reg, col_reg}<16'b0111100000101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111100000101110) && ({row_reg, col_reg}<16'b0111100000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100000110001) && ({row_reg, col_reg}<16'b0111100000110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111100000110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111100000110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111100000110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111100000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111100000110111) && ({row_reg, col_reg}<16'b0111100000111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111100000111001) && ({row_reg, col_reg}<16'b0111100000111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111100000111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111100000111101) && ({row_reg, col_reg}<16'b0111100000111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111100000111111) && ({row_reg, col_reg}<16'b0111100001000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111100001000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111100001000100) && ({row_reg, col_reg}<16'b0111100001000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111100001000111) && ({row_reg, col_reg}<16'b0111100001001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111100001001001) && ({row_reg, col_reg}<16'b0111100001001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111100001001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111100001001101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0111100001001110) && ({row_reg, col_reg}<16'b0111100001010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111100001010000) && ({row_reg, col_reg}<16'b0111100001010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111100001010011) && ({row_reg, col_reg}<16'b0111100001010101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111100001010101) && ({row_reg, col_reg}<16'b0111100001011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111100001011000) && ({row_reg, col_reg}<16'b0111100001011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0111100001011010) && ({row_reg, col_reg}<16'b0111100001011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111100001011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111100001011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111100001011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111100001011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111100001100000) && ({row_reg, col_reg}<16'b0111100001100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111100001100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111100001100011) && ({row_reg, col_reg}<16'b0111100001100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111100001100110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111100001100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111100001101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111100001101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111100001101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111100001101011) && ({row_reg, col_reg}<16'b0111100001110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111100001110001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111100001110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111100001110011) && ({row_reg, col_reg}<16'b0111100001110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111100001110101) && ({row_reg, col_reg}<16'b0111100001110111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111100001110111) && ({row_reg, col_reg}<16'b0111100001111100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111100001111100) && ({row_reg, col_reg}<16'b0111100010000100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111100010000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111100010000101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111100010000110) && ({row_reg, col_reg}<16'b0111100010010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111100010010000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111100010010001)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0111100010010010) && ({row_reg, col_reg}<16'b0111100010010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111100010010100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111100010010101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0111100010010110) && ({row_reg, col_reg}<16'b0111100010011000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0111100010011000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0111100010011001) && ({row_reg, col_reg}<16'b0111100010011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111100010011100) && ({row_reg, col_reg}<16'b0111100010100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111100010100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111100010100010) && ({row_reg, col_reg}<16'b0111100010101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111100010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111100010101001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111100010101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111100010101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111100010101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111100010101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111100010101110) && ({row_reg, col_reg}<16'b0111100010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111100010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111100010110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111100010110101) && ({row_reg, col_reg}<16'b0111100010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100010111100) && ({row_reg, col_reg}<16'b0111100010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100010111110) && ({row_reg, col_reg}<16'b0111100011000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111100011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100011000001) && ({row_reg, col_reg}<16'b0111100011000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111100011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111100011000110) && ({row_reg, col_reg}<16'b0111100011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100011010001) && ({row_reg, col_reg}<16'b0111100011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111100011110000) && ({row_reg, col_reg}<16'b0111100011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111100011110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111100011110011) && ({row_reg, col_reg}<16'b0111100011110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111100011110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111100011111000) && ({row_reg, col_reg}<16'b0111100011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111100011111011)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0111100011111100) && ({row_reg, col_reg}<16'b0111100100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111100100000000) && ({row_reg, col_reg}<16'b0111100100000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100100000100) && ({row_reg, col_reg}<16'b0111100100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100100001101) && ({row_reg, col_reg}<16'b0111100100001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111100100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111100100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111100100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111100100010010) && ({row_reg, col_reg}<16'b0111100100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111100100100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100100100110) && ({row_reg, col_reg}<16'b0111100100101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111100100101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100100101011) && ({row_reg, col_reg}<16'b0111100100101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111100100101110) && ({row_reg, col_reg}<16'b0111100100110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100100110010) && ({row_reg, col_reg}<16'b0111100100110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100100110100) && ({row_reg, col_reg}<16'b0111100100110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111100100110111) && ({row_reg, col_reg}<16'b0111100100111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111100100111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111100100111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100100111011) && ({row_reg, col_reg}<16'b0111100100111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111100100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100100111111) && ({row_reg, col_reg}<16'b0111100101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100101000001) && ({row_reg, col_reg}<16'b0111100101001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111100101001101) && ({row_reg, col_reg}<16'b0111100101011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111100101011010) && ({row_reg, col_reg}<16'b0111100101011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111100101011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111100101011101) && ({row_reg, col_reg}<16'b0111100101011111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111100101011111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0111100101100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111100101100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111100101100010) && ({row_reg, col_reg}<16'b0111100101100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111100101100110) && ({row_reg, col_reg}<16'b0111100101101000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111100101101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111100101101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111100101101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111100101101011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111100101101100) && ({row_reg, col_reg}<16'b0111100101101110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111100101101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111100101101111) && ({row_reg, col_reg}<16'b0111100101110001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111100101110001) && ({row_reg, col_reg}<16'b0111100101111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111100101111001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111100101111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111100101111011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111100101111100) && ({row_reg, col_reg}<16'b0111100110001000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111100110001000) && ({row_reg, col_reg}<16'b0111100110001100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111100110001100) && ({row_reg, col_reg}<16'b0111100110001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111100110001111) && ({row_reg, col_reg}<16'b0111100110010001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111100110010001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111100110010010)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0111100110010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111100110010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111100110010101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111100110010110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0111100110010111)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0111100110011000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0111100110011001) && ({row_reg, col_reg}<16'b0111100110011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111100110011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111100110011111) && ({row_reg, col_reg}<16'b0111100110101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111100110101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111100110101010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0111100110101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111100110101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111100110101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111100110101110) && ({row_reg, col_reg}<16'b0111100110110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111100110110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111100110110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111100110110010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0111100110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111100110110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111100110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100110110110) && ({row_reg, col_reg}<16'b0111100110111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111100110111001) && ({row_reg, col_reg}<16'b0111100110111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100110111100) && ({row_reg, col_reg}<16'b0111100110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100110111110) && ({row_reg, col_reg}<16'b0111100111000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111100111000000) && ({row_reg, col_reg}<16'b0111100111000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111100111000100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111100111000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111100111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111100111000111) && ({row_reg, col_reg}<16'b0111100111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100111010001) && ({row_reg, col_reg}<16'b0111100111110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111100111110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111100111110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100111110010) && ({row_reg, col_reg}<16'b0111100111110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111100111110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100111110111) && ({row_reg, col_reg}<16'b0111100111111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100111111100) && ({row_reg, col_reg}<16'b0111100111111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111100111111110)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}==16'b0111100111111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111101000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101000000001) && ({row_reg, col_reg}<16'b0111101000000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101000000101) && ({row_reg, col_reg}<16'b0111101000001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101000001000) && ({row_reg, col_reg}<16'b0111101000001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101000001010) && ({row_reg, col_reg}<16'b0111101000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101000001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111101000001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111101000001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111101000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101000010010) && ({row_reg, col_reg}<16'b0111101000100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111101000100100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111101000100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101000100110) && ({row_reg, col_reg}<16'b0111101000101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111101000101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101000101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111101000101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111101000101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101000101110) && ({row_reg, col_reg}<16'b0111101000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101000110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101000110010) && ({row_reg, col_reg}<16'b0111101000110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111101000110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111101000110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111101000110110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0111101000110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111101000111001) && ({row_reg, col_reg}<16'b0111101000111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101000111100) && ({row_reg, col_reg}<16'b0111101000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111101000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101000111111) && ({row_reg, col_reg}<16'b0111101001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101001000001) && ({row_reg, col_reg}<16'b0111101001000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111101001000011) && ({row_reg, col_reg}<16'b0111101001011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101001011011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0111101001011100) && ({row_reg, col_reg}<16'b0111101001011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111101001011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111101001011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0111101001100000) && ({row_reg, col_reg}<16'b0111101001100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111101001100011) && ({row_reg, col_reg}<16'b0111101001100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111101001100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111101001100110) && ({row_reg, col_reg}<16'b0111101001101000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111101001101000) && ({row_reg, col_reg}<16'b0111101001101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101001101010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111101001101011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111101001101100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111101001101101) && ({row_reg, col_reg}<16'b0111101001101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0111101001101111) && ({row_reg, col_reg}<16'b0111101001110010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111101001110010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111101001110011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111101001110100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111101001110101) && ({row_reg, col_reg}<16'b0111101001111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111101001111110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111101001111111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111101010000000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111101010000001) && ({row_reg, col_reg}<16'b0111101010000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111101010000111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111101010001000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111101010001001) && ({row_reg, col_reg}<16'b0111101010001100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111101010001100) && ({row_reg, col_reg}<16'b0111101010001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111101010001110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111101010001111) && ({row_reg, col_reg}<16'b0111101010010001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111101010010001) && ({row_reg, col_reg}<16'b0111101010010011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111101010010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111101010010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0111101010010101) && ({row_reg, col_reg}<16'b0111101010011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111101010011001) && ({row_reg, col_reg}<16'b0111101010011011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111101010011011) && ({row_reg, col_reg}<16'b0111101010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101010100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111101010101000) && ({row_reg, col_reg}<16'b0111101010101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101010101100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0111101010101101) && ({row_reg, col_reg}<16'b0111101010101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101010101111) && ({row_reg, col_reg}<16'b0111101010110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111101010110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111101010110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111101010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111101010110101) && ({row_reg, col_reg}<16'b0111101010110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111101010110111) && ({row_reg, col_reg}<16'b0111101010111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111101010111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111101010111010) && ({row_reg, col_reg}<16'b0111101010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111101010111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101010111101) && ({row_reg, col_reg}<16'b0111101011000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111101011000000) && ({row_reg, col_reg}<16'b0111101011000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101011000100) && ({row_reg, col_reg}<16'b0111101011001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101011001000) && ({row_reg, col_reg}<16'b0111101011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101011001010) && ({row_reg, col_reg}<16'b0111101011001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101011001100) && ({row_reg, col_reg}<16'b0111101011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101011010001) && ({row_reg, col_reg}<16'b0111101011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111101011110000) && ({row_reg, col_reg}<16'b0111101011110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101011110010) && ({row_reg, col_reg}<16'b0111101011110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111101011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111101011110110) && ({row_reg, col_reg}<16'b0111101011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111101011111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101011111100) && ({row_reg, col_reg}<16'b0111101011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111101011111110)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}==16'b0111101011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111101100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101100000001) && ({row_reg, col_reg}<16'b0111101100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101100000101) && ({row_reg, col_reg}<16'b0111101100001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101100001001) && ({row_reg, col_reg}<16'b0111101100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101100001011) && ({row_reg, col_reg}<16'b0111101100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101100001101) && ({row_reg, col_reg}<16'b0111101100010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111101100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101100010010) && ({row_reg, col_reg}<16'b0111101100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111101100100101) && ({row_reg, col_reg}<16'b0111101100101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111101100101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101100101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111101100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111101100101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101100101110) && ({row_reg, col_reg}<16'b0111101100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101100110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111101100110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111101100110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111101100110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111101100110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111101100110110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0111101100110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101100111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111101100111001) && ({row_reg, col_reg}<16'b0111101100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111101100111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101100111100) && ({row_reg, col_reg}<16'b0111101100111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111101100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101100111111) && ({row_reg, col_reg}<16'b0111101101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111101101000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111101101000010) && ({row_reg, col_reg}<16'b0111101101000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101101000100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111101101000101) && ({row_reg, col_reg}<16'b0111101101001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111101101001110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111101101001111) && ({row_reg, col_reg}<16'b0111101101011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101101011011) && ({row_reg, col_reg}<16'b0111101101011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111101101011110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111101101011111)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0111101101100000) && ({row_reg, col_reg}<16'b0111101101101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111101101101000) && ({row_reg, col_reg}<16'b0111101101101010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111101101101010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111101101101011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111101101101100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111101101101101) && ({row_reg, col_reg}<16'b0111101101110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111101101110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111101101110001) && ({row_reg, col_reg}<16'b0111101101110100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111101101110100) && ({row_reg, col_reg}<16'b0111101101110111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111101101110111) && ({row_reg, col_reg}<16'b0111101101111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111101101111100) && ({row_reg, col_reg}<16'b0111101101111110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111101101111110) && ({row_reg, col_reg}<16'b0111101110000001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0111101110000001) && ({row_reg, col_reg}<16'b0111101110000111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111101110000111) && ({row_reg, col_reg}<16'b0111101110001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111101110001100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111101110001101) && ({row_reg, col_reg}<16'b0111101110001111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111101110001111) && ({row_reg, col_reg}<16'b0111101110010001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111101110010001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111101110010010) && ({row_reg, col_reg}<16'b0111101110010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111101110010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101110010101) && ({row_reg, col_reg}<16'b0111101110010111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0111101110010111) && ({row_reg, col_reg}<16'b0111101110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101110100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111101110101000) && ({row_reg, col_reg}<16'b0111101110101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101110101100) && ({row_reg, col_reg}<16'b0111101110110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111101110110001) && ({row_reg, col_reg}<16'b0111101110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101110110011) && ({row_reg, col_reg}<16'b0111101110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111101110110101) && ({row_reg, col_reg}<16'b0111101110110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111101110110111) && ({row_reg, col_reg}<16'b0111101110111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111101110111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111101110111010) && ({row_reg, col_reg}<16'b0111101110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101110111101) && ({row_reg, col_reg}<16'b0111101110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111101110111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111101111000000) && ({row_reg, col_reg}<16'b0111101111000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101111000010) && ({row_reg, col_reg}<16'b0111101111000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101111000111) && ({row_reg, col_reg}<16'b0111101111001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101111001010) && ({row_reg, col_reg}<16'b0111101111001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101111001100) && ({row_reg, col_reg}<16'b0111101111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101111010001) && ({row_reg, col_reg}<16'b0111101111101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111101111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101111110000) && ({row_reg, col_reg}<16'b0111101111110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101111110010) && ({row_reg, col_reg}<16'b0111101111110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111101111110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101111110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111101111110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111101111110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101111111000) && ({row_reg, col_reg}<16'b0111101111111011)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0111101111111011) && ({row_reg, col_reg}<16'b0111110000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111110000000000) && ({row_reg, col_reg}<16'b0111110000000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110000000100) && ({row_reg, col_reg}<16'b0111110000001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110000001001) && ({row_reg, col_reg}<16'b0111110000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111110000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110000001101) && ({row_reg, col_reg}<16'b0111110000001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110000001111) && ({row_reg, col_reg}<16'b0111110000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110000010010) && ({row_reg, col_reg}<16'b0111110000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111110000100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110000100110) && ({row_reg, col_reg}<16'b0111110000101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110000101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111110000101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111110000101101) && ({row_reg, col_reg}<16'b0111110000101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110000101111) && ({row_reg, col_reg}<16'b0111110000110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110000110001) && ({row_reg, col_reg}<16'b0111110000110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111110000110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110000110100) && ({row_reg, col_reg}<16'b0111110000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111110000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111110000110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111110000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110000111001) && ({row_reg, col_reg}<16'b0111110000111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110000111100) && ({row_reg, col_reg}<16'b0111110000111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111110000111111) && ({row_reg, col_reg}<16'b0111110001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111110001000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111110001000010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0111110001000011) && ({row_reg, col_reg}<16'b0111110001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110001000101) && ({row_reg, col_reg}<16'b0111110001001001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111110001001001) && ({row_reg, col_reg}<16'b0111110001001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111110001001111) && ({row_reg, col_reg}<16'b0111110001010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111110001010010) && ({row_reg, col_reg}<16'b0111110001010101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111110001010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111110001010110) && ({row_reg, col_reg}<16'b0111110001011000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111110001011000) && ({row_reg, col_reg}<16'b0111110001011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110001011110) && ({row_reg, col_reg}<16'b0111110001100000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111110001100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111110001100001) && ({row_reg, col_reg}<16'b0111110001100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111110001100101) && ({row_reg, col_reg}<16'b0111110001100111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111110001100111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111110001101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111110001101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111110001101010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0111110001101011) && ({row_reg, col_reg}<16'b0111110001101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111110001101101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111110001101110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111110001101111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111110001110000) && ({row_reg, col_reg}<16'b0111110001110011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111110001110011) && ({row_reg, col_reg}<16'b0111110001110110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111110001110110) && ({row_reg, col_reg}<16'b0111110001111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111110001111000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111110001111001) && ({row_reg, col_reg}<16'b0111110001111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111110001111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111110001111100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111110001111101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111110001111110) && ({row_reg, col_reg}<16'b0111110010000001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0111110010000001) && ({row_reg, col_reg}<16'b0111110010000101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111110010000101) && ({row_reg, col_reg}<16'b0111110010000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111110010000111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111110010001000) && ({row_reg, col_reg}<16'b0111110010001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111110010001101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111110010001110) && ({row_reg, col_reg}<16'b0111110010010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111110010010010) && ({row_reg, col_reg}<16'b0111110010010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111110010010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110010010101) && ({row_reg, col_reg}<16'b0111110010011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111110010011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110010011010) && ({row_reg, col_reg}<16'b0111110010011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110010011100) && ({row_reg, col_reg}<16'b0111110010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110010100011) && ({row_reg, col_reg}<16'b0111110010101010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111110010101010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111110010101011) && ({row_reg, col_reg}<16'b0111110010101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111110010101111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111110010110000) && ({row_reg, col_reg}<16'b0111110010110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111110010110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111110010110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111110010110100) && ({row_reg, col_reg}<16'b0111110010110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111110010110111) && ({row_reg, col_reg}<16'b0111110010111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110010111001) && ({row_reg, col_reg}<16'b0111110010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110010111101) && ({row_reg, col_reg}<16'b0111110010111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111110010111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111110011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110011000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110011000010) && ({row_reg, col_reg}<16'b0111110011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111110011000100) && ({row_reg, col_reg}<16'b0111110011000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110011000111) && ({row_reg, col_reg}<16'b0111110011001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110011001011) && ({row_reg, col_reg}<16'b0111110011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111110011001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111110011001111) && ({row_reg, col_reg}<16'b0111110011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110011010001) && ({row_reg, col_reg}<16'b0111110011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111110011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110011110000) && ({row_reg, col_reg}<16'b0111110011110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110011110010) && ({row_reg, col_reg}<16'b0111110011110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110011110110) && ({row_reg, col_reg}<16'b0111110011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111110011111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111110011111010)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0111110011111011) && ({row_reg, col_reg}<16'b0111110100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111110100000000) && ({row_reg, col_reg}<16'b0111110100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110100000010) && ({row_reg, col_reg}<16'b0111110100001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110100001000) && ({row_reg, col_reg}<16'b0111110100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110100001011) && ({row_reg, col_reg}<16'b0111110100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110100001101) && ({row_reg, col_reg}<16'b0111110100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110100001111) && ({row_reg, col_reg}<16'b0111110100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111110100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110100010010) && ({row_reg, col_reg}<16'b0111110100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111110100100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110100100110) && ({row_reg, col_reg}<16'b0111110100101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110100101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111110100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111110100101101) && ({row_reg, col_reg}<16'b0111110100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110100110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111110100110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111110100110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111110100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111110100110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111110100110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111110100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111110100110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111110100111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110100111001) && ({row_reg, col_reg}<16'b0111110100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111110100111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110100111100) && ({row_reg, col_reg}<16'b0111110100111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111110100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110100111111) && ({row_reg, col_reg}<16'b0111110101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111110101000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111110101000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111110101000011) && ({row_reg, col_reg}<16'b0111110101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110101000110) && ({row_reg, col_reg}<16'b0111110101001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110101001011) && ({row_reg, col_reg}<16'b0111110101010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111110101010010) && ({row_reg, col_reg}<16'b0111110101011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111110101011001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111110101011010) && ({row_reg, col_reg}<16'b0111110101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111110101011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111110101011111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0111110101100000) && ({row_reg, col_reg}<16'b0111110101100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111110101100110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111110101100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111110101101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111110101101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111110101101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110101101011) && ({row_reg, col_reg}<16'b0111110101101101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111110101101101) && ({row_reg, col_reg}<16'b0111110101110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111110101110011) && ({row_reg, col_reg}<16'b0111110101110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111110101110101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111110101110110) && ({row_reg, col_reg}<16'b0111110101111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111110101111000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111110101111001) && ({row_reg, col_reg}<16'b0111110101111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111110101111100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111110101111101) && ({row_reg, col_reg}<16'b0111110101111111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111110101111111) && ({row_reg, col_reg}<16'b0111110110000001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111110110000001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111110110000010) && ({row_reg, col_reg}<16'b0111110110000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111110110000100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111110110000101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111110110000110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111110110000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111110110001000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111110110001001) && ({row_reg, col_reg}<16'b0111110110001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111110110001111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111110110010000) && ({row_reg, col_reg}<16'b0111110110010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110110010101) && ({row_reg, col_reg}<16'b0111110110011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110110011000) && ({row_reg, col_reg}<16'b0111110110011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111110110011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111110110011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111110110011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111110110100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111110110100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111110110100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110110100011) && ({row_reg, col_reg}<16'b0111110110101110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111110110101110) && ({row_reg, col_reg}<16'b0111110110110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110110110000) && ({row_reg, col_reg}<16'b0111110110110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110110110010) && ({row_reg, col_reg}<16'b0111110110110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111110110110101) && ({row_reg, col_reg}<16'b0111110110111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111110110111001) && ({row_reg, col_reg}<16'b0111110111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111110111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110111000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110111000010) && ({row_reg, col_reg}<16'b0111110111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111110111000100) && ({row_reg, col_reg}<16'b0111110111001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111110111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110111001001) && ({row_reg, col_reg}<16'b0111110111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110111001011) && ({row_reg, col_reg}<16'b0111110111001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110111001101) && ({row_reg, col_reg}<16'b0111110111001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111110111001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111110111010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110111010001) && ({row_reg, col_reg}<16'b0111110111110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111110111110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110111110001) && ({row_reg, col_reg}<16'b0111110111110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110111110011) && ({row_reg, col_reg}<16'b0111110111110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110111110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111110111110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111110111110111) && ({row_reg, col_reg}<16'b0111110111111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111110111111010)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0111110111111011) && ({row_reg, col_reg}<16'b0111111000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111111000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111000000001) && ({row_reg, col_reg}<16'b0111111000001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111000001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111000001011) && ({row_reg, col_reg}<16'b0111111000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111000001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111000001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111111000001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111000010000) && ({row_reg, col_reg}<16'b0111111000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111000010010) && ({row_reg, col_reg}<16'b0111111000100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111111000100100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111111000100101) && ({row_reg, col_reg}<16'b0111111000101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111000101010) && ({row_reg, col_reg}<16'b0111111000101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111000101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111111000101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111111000101110) && ({row_reg, col_reg}<16'b0111111000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111000110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111000110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111111000110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111000110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111111000110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111111000110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111111000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111111000110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111111000111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111111000111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111111000111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111111000111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111000111101) && ({row_reg, col_reg}<16'b0111111000111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111111000111111) && ({row_reg, col_reg}<16'b0111111001000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111111001000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111111001000010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0111111001000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111001000100) && ({row_reg, col_reg}<16'b0111111001001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111111001001000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0111111001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111001001010) && ({row_reg, col_reg}<16'b0111111001010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111001010001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111111001010010) && ({row_reg, col_reg}<16'b0111111001011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111111001011010) && ({row_reg, col_reg}<16'b0111111001011101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111111001011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111111001011110) && ({row_reg, col_reg}<16'b0111111001100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111001100000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111111001100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111111001100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111111001100011) && ({row_reg, col_reg}<16'b0111111001100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111001100101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111111001100110) && ({row_reg, col_reg}<16'b0111111001101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111111001101000) && ({row_reg, col_reg}<16'b0111111001110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111001110000) && ({row_reg, col_reg}<16'b0111111001110010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111111001110010) && ({row_reg, col_reg}<16'b0111111001110100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111111001110100) && ({row_reg, col_reg}<16'b0111111001110110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111111001110110) && ({row_reg, col_reg}<16'b0111111001111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0111111001111000) && ({row_reg, col_reg}<16'b0111111001111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111111001111011) && ({row_reg, col_reg}<16'b0111111001111110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111111001111110) && ({row_reg, col_reg}<16'b0111111010000000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111111010000000) && ({row_reg, col_reg}<16'b0111111010000010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111111010000010) && ({row_reg, col_reg}<16'b0111111010000100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111111010000100) && ({row_reg, col_reg}<16'b0111111010000110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111111010000110) && ({row_reg, col_reg}<16'b0111111010001001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111111010001001) && ({row_reg, col_reg}<16'b0111111010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111111010001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111111010001101) && ({row_reg, col_reg}<16'b0111111010011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111010011101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111111010011110) && ({row_reg, col_reg}<16'b0111111010100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111111010100100) && ({row_reg, col_reg}<16'b0111111010100110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111111010100110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111111010100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111111010101000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111111010101001) && ({row_reg, col_reg}<16'b0111111010101110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111010101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111010101111) && ({row_reg, col_reg}<16'b0111111010110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111111010110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111010110010) && ({row_reg, col_reg}<16'b0111111010110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111111010110110) && ({row_reg, col_reg}<16'b0111111010111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111010111011) && ({row_reg, col_reg}<16'b0111111011000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111111011000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111111011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111011000010) && ({row_reg, col_reg}<16'b0111111011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111111011000100) && ({row_reg, col_reg}<16'b0111111011001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111011001001) && ({row_reg, col_reg}<16'b0111111011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111011001011) && ({row_reg, col_reg}<16'b0111111011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111011001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111111011001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111011010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111011010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111111011010010) && ({row_reg, col_reg}<16'b0111111011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111111011101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111011110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111011110001) && ({row_reg, col_reg}<16'b0111111011110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111011110011) && ({row_reg, col_reg}<16'b0111111011110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111011110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111111011110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111011111000) && ({row_reg, col_reg}<16'b0111111011111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111011111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111011111011) && ({row_reg, col_reg}<16'b0111111011111111)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}==16'b0111111011111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111100000001) && ({row_reg, col_reg}<16'b0111111100001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111100001011) && ({row_reg, col_reg}<16'b0111111100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111100001101) && ({row_reg, col_reg}<16'b0111111100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111111100001111) && ({row_reg, col_reg}<16'b0111111100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111111100010011) && ({row_reg, col_reg}<16'b0111111100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111111100100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111111100100110) && ({row_reg, col_reg}<16'b0111111100101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111100101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111111100101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111111100101110) && ({row_reg, col_reg}<16'b0111111100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111100110000) && ({row_reg, col_reg}<16'b0111111100110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111100110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111111100110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111111100110101) && ({row_reg, col_reg}<16'b0111111100110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111100110111) && ({row_reg, col_reg}<16'b0111111100111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111100111001) && ({row_reg, col_reg}<16'b0111111100111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111100111100) && ({row_reg, col_reg}<16'b0111111100111110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111100111110) && ({row_reg, col_reg}<16'b0111111101000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111111101000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111101000101) && ({row_reg, col_reg}<16'b0111111101001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111111101001010) && ({row_reg, col_reg}<16'b0111111101001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111101001101) && ({row_reg, col_reg}<16'b0111111101010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111101010010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111111101010011) && ({row_reg, col_reg}<16'b0111111101011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111111101011110) && ({row_reg, col_reg}<16'b0111111101101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111101101011) && ({row_reg, col_reg}<16'b0111111101101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111101101101) && ({row_reg, col_reg}<16'b0111111101110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111101110011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111111101110100) && ({row_reg, col_reg}<16'b0111111101111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111111101111010) && ({row_reg, col_reg}<16'b0111111110000101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111111110000101) && ({row_reg, col_reg}<16'b0111111110001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111111110001001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111111110001010) && ({row_reg, col_reg}<16'b0111111110001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111110001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111110001111) && ({row_reg, col_reg}<16'b0111111110010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111110010110) && ({row_reg, col_reg}<16'b0111111110011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111111110011001) && ({row_reg, col_reg}<16'b0111111110011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111111110011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111110011101) && ({row_reg, col_reg}<16'b0111111110100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111111110100100) && ({row_reg, col_reg}<16'b0111111110100110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111111110100110) && ({row_reg, col_reg}<16'b0111111110101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111111110101000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111111110101001) && ({row_reg, col_reg}<16'b0111111110101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111110101100) && ({row_reg, col_reg}<16'b0111111110101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111110101110) && ({row_reg, col_reg}<16'b0111111110110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111111110110001) && ({row_reg, col_reg}<16'b0111111110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111111110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111111110111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111111110111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111110111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111111110111100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0111111110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111110111110) && ({row_reg, col_reg}<16'b0111111111000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111111000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111111111000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111111111000100) && ({row_reg, col_reg}<16'b0111111111001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111111001001) && ({row_reg, col_reg}<16'b0111111111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111111111001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111111001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111111001101) && ({row_reg, col_reg}<16'b0111111111010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111111010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111111010001) && ({row_reg, col_reg}<16'b0111111111101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111111111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111111110000) && ({row_reg, col_reg}<16'b0111111111110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111111110011) && ({row_reg, col_reg}<16'b0111111111110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111111110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111111111110110) && ({row_reg, col_reg}<16'b0111111111111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111111111111000) && ({row_reg, col_reg}<16'b0111111111111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111111111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111111111011) && ({row_reg, col_reg}<16'b0111111111111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0111111111111110) && ({row_reg, col_reg}<16'b1000000000000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000000000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000000000001) && ({row_reg, col_reg}<16'b1000000000001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000000001001) && ({row_reg, col_reg}<16'b1000000000001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000000001011) && ({row_reg, col_reg}<16'b1000000000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000000000010011) && ({row_reg, col_reg}<16'b1000000000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000000000100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000000000100110) && ({row_reg, col_reg}<16'b1000000000101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000000101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000000000101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000000000101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000000000101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000000000101110) && ({row_reg, col_reg}<16'b1000000000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000000110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000000000110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000000110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000000110100) && ({row_reg, col_reg}<16'b1000000000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000000000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000000110111) && ({row_reg, col_reg}<16'b1000000000111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000000111111) && ({row_reg, col_reg}<16'b1000000001000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000000001000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000001000100) && ({row_reg, col_reg}<16'b1000000001000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000001000111) && ({row_reg, col_reg}<16'b1000000001001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000000001001101) && ({row_reg, col_reg}<16'b1000000001010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000001010000) && ({row_reg, col_reg}<16'b1000000001010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000001010011) && ({row_reg, col_reg}<16'b1000000001011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000000001011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000000001011111) && ({row_reg, col_reg}<16'b1000000001111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000000001111000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000000001111001) && ({row_reg, col_reg}<16'b1000000001111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000000001111101) && ({row_reg, col_reg}<16'b1000000010000000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b1000000010000000) && ({row_reg, col_reg}<16'b1000000010000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000000010000101) && ({row_reg, col_reg}<16'b1000000010000111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000000010000111) && ({row_reg, col_reg}<16'b1000000010001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000000010001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000010001111) && ({row_reg, col_reg}<16'b1000000010010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000010010010) && ({row_reg, col_reg}<16'b1000000010010100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000000010010100) && ({row_reg, col_reg}<16'b1000000010010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000000010010110) && ({row_reg, col_reg}<16'b1000000010011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000000010011011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000000010011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000010011101) && ({row_reg, col_reg}<16'b1000000010100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000000010100101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000000010100110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000000010100111) && ({row_reg, col_reg}<16'b1000000010101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000000010101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000010101100) && ({row_reg, col_reg}<16'b1000000010101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000000010101110) && ({row_reg, col_reg}<16'b1000000010110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000010110010) && ({row_reg, col_reg}<16'b1000000010110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000010110100) && ({row_reg, col_reg}<16'b1000000010111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000010111001) && ({row_reg, col_reg}<16'b1000000010111100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000000010111100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000000010111101) && ({row_reg, col_reg}<16'b1000000011000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000000011000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000000011000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000000011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000000011000100) && ({row_reg, col_reg}<16'b1000000011001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000000011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000011001001) && ({row_reg, col_reg}<16'b1000000011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000000011001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000000011001100) && ({row_reg, col_reg}<16'b1000000011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000000011001111) && ({row_reg, col_reg}<16'b1000000011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000011010001) && ({row_reg, col_reg}<16'b1000000011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000000011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000011110000) && ({row_reg, col_reg}<16'b1000000011110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000011110011) && ({row_reg, col_reg}<16'b1000000011110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000011110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000000011110110) && ({row_reg, col_reg}<16'b1000000011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000000011111001) && ({row_reg, col_reg}<16'b1000000011111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000000011111011) && ({row_reg, col_reg}<16'b1000000011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000000011111110)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}==16'b1000000011111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000100000001) && ({row_reg, col_reg}<16'b1000000100001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000100001001) && ({row_reg, col_reg}<16'b1000000100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000100001100) && ({row_reg, col_reg}<16'b1000000100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000100010010) && ({row_reg, col_reg}<16'b1000000100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000000100100110) && ({row_reg, col_reg}<16'b1000000100101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000100101001) && ({row_reg, col_reg}<16'b1000000100101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000000100101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000000100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000000100101101) && ({row_reg, col_reg}<16'b1000000100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000100110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000100110101) && ({row_reg, col_reg}<16'b1000000100110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000000100110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000100111000) && ({row_reg, col_reg}<16'b1000000100111110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000100111110) && ({row_reg, col_reg}<16'b1000000101000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000000101000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1000000101000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000101000010) && ({row_reg, col_reg}<16'b1000000101000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000101000111) && ({row_reg, col_reg}<16'b1000000101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000000101001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000000101001010) && ({row_reg, col_reg}<16'b1000000101001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000000101001101) && ({row_reg, col_reg}<16'b1000000101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000000101001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000000101010000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1000000101010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000101010010) && ({row_reg, col_reg}<16'b1000000101010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000101010101) && ({row_reg, col_reg}<16'b1000000101011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000000101011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000000101011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000101100000) && ({row_reg, col_reg}<16'b1000000101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000101100010) && ({row_reg, col_reg}<16'b1000000101100100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000101100100) && ({row_reg, col_reg}<16'b1000000101100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000000101100111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000000101101000) && ({row_reg, col_reg}<16'b1000000101101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000101101011) && ({row_reg, col_reg}<16'b1000000101101110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000000101101110) && ({row_reg, col_reg}<16'b1000000101110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000000101110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000101110111) && ({row_reg, col_reg}<16'b1000000101111100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000000101111100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000000101111101) && ({row_reg, col_reg}<16'b1000000110000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000000110000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000000110000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000000110000011) && ({row_reg, col_reg}<16'b1000000110010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000110010001) && ({row_reg, col_reg}<16'b1000000110011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000000110011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000000110011101) && ({row_reg, col_reg}<16'b1000000110100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000000110100100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000000110100101) && ({row_reg, col_reg}<16'b1000000110101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000110101000) && ({row_reg, col_reg}<16'b1000000110101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000000110101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000000110101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000000110101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000110101110) && ({row_reg, col_reg}<16'b1000000110111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000110111000) && ({row_reg, col_reg}<16'b1000000110111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000110111100) && ({row_reg, col_reg}<16'b1000000110111110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000110111110) && ({row_reg, col_reg}<16'b1000000111000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000000111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000111000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000000111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000000111000100) && ({row_reg, col_reg}<16'b1000000111001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000000111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000111001001) && ({row_reg, col_reg}<16'b1000000111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000111001011) && ({row_reg, col_reg}<16'b1000000111001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000000111001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000000111001111) && ({row_reg, col_reg}<16'b1000000111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000111010001) && ({row_reg, col_reg}<16'b1000000111101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000000111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000111110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000000111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000111110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000000111110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000000111110100) && ({row_reg, col_reg}<16'b1000000111110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000111110110) && ({row_reg, col_reg}<16'b1000000111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000000111111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000000111111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000111111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000000111111100) && ({row_reg, col_reg}<16'b1000000111111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000000111111110)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}==16'b1000000111111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001000000001) && ({row_reg, col_reg}<16'b1000001000001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001000001010) && ({row_reg, col_reg}<16'b1000001000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001000001100) && ({row_reg, col_reg}<16'b1000001000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000001000010010) && ({row_reg, col_reg}<16'b1000001000100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000001000100110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000001000100111) && ({row_reg, col_reg}<16'b1000001000101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001000101011) && ({row_reg, col_reg}<16'b1000001000101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000001000101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000001000101110) && ({row_reg, col_reg}<16'b1000001000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001000110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000001000110010) && ({row_reg, col_reg}<16'b1000001000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001000110101) && ({row_reg, col_reg}<16'b1000001000111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000001000111001) && ({row_reg, col_reg}<16'b1000001000111100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001000111100) && ({row_reg, col_reg}<16'b1000001001000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001001000001) && ({row_reg, col_reg}<16'b1000001001000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001001000111) && ({row_reg, col_reg}<16'b1000001001001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000001001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001001001011) && ({row_reg, col_reg}<16'b1000001001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001001001111) && ({row_reg, col_reg}<16'b1000001001010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000001001010001) && ({row_reg, col_reg}<16'b1000001001010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001001010011) && ({row_reg, col_reg}<16'b1000001001010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000001001010111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000001001011000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000001001011001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000001001011010) && ({row_reg, col_reg}<16'b1000001001011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000001001011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000001001011110) && ({row_reg, col_reg}<16'b1000001001100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001001100000) && ({row_reg, col_reg}<16'b1000001001100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001001100010) && ({row_reg, col_reg}<16'b1000001001100100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001001100100) && ({row_reg, col_reg}<16'b1000001001101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000001001101111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000001001110000) && ({row_reg, col_reg}<16'b1000001001110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001001110111) && ({row_reg, col_reg}<16'b1000001001111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001001111001) && ({row_reg, col_reg}<16'b1000001010001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001010001101) && ({row_reg, col_reg}<16'b1000001010100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000001010100011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000001010100100) && ({row_reg, col_reg}<16'b1000001010100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001010100110) && ({row_reg, col_reg}<16'b1000001010101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001010101101) && ({row_reg, col_reg}<16'b1000001010111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001010111000) && ({row_reg, col_reg}<16'b1000001010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000001010111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000001010111011) && ({row_reg, col_reg}<16'b1000001010111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000001010111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000001011000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000001011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001011000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000001011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000001011000100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000001011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000001011000110) && ({row_reg, col_reg}<16'b1000001011001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000001011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001011001001) && ({row_reg, col_reg}<16'b1000001011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000001011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000001011001100) && ({row_reg, col_reg}<16'b1000001011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000001011001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000001011001111) && ({row_reg, col_reg}<16'b1000001011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001011010001) && ({row_reg, col_reg}<16'b1000001011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000001011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000001011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001011110010) && ({row_reg, col_reg}<16'b1000001011110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000001011110100) && ({row_reg, col_reg}<16'b1000001011110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001011110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000001011110111) && ({row_reg, col_reg}<16'b1000001011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000001011111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000001011111010) && ({row_reg, col_reg}<16'b1000001011111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001011111100) && ({row_reg, col_reg}<16'b1000001011111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b1000001011111110) && ({row_reg, col_reg}<16'b1000001100000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000001100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001100000001) && ({row_reg, col_reg}<16'b1000001100001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001100001010) && ({row_reg, col_reg}<16'b1000001100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001100001100) && ({row_reg, col_reg}<16'b1000001100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001100001111) && ({row_reg, col_reg}<16'b1000001100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000001100010010) && ({row_reg, col_reg}<16'b1000001100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000001100100110) && ({row_reg, col_reg}<16'b1000001100101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001100101001) && ({row_reg, col_reg}<16'b1000001100101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001100101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000001100101101) && ({row_reg, col_reg}<16'b1000001100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001100110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000001100110110) && ({row_reg, col_reg}<16'b1000001100111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001100111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000001100111010) && ({row_reg, col_reg}<16'b1000001100111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001100111101) && ({row_reg, col_reg}<16'b1000001100111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000001100111111) && ({row_reg, col_reg}<16'b1000001101000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001101000111) && ({row_reg, col_reg}<16'b1000001101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001101001001) && ({row_reg, col_reg}<16'b1000001101001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000001101001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001101001111) && ({row_reg, col_reg}<16'b1000001101010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000001101010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000001101010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001101010011) && ({row_reg, col_reg}<16'b1000001101010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000001101010101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1000001101010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001101010111) && ({row_reg, col_reg}<16'b1000001101011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001101011011) && ({row_reg, col_reg}<16'b1000001101011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000001101011101) && ({row_reg, col_reg}<16'b1000001101011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001101011111) && ({row_reg, col_reg}<16'b1000001101100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000001101100001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1000001101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000001101100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000001101100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000001101100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b1000001101100110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b1000001101100111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b1000001101101000) && ({row_reg, col_reg}<16'b1000001101101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000001101101111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000001101110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000001101110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000001101110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000001101110011) && ({row_reg, col_reg}<16'b1000001101110101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000001101110101) && ({row_reg, col_reg}<16'b1000001110001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000001110001000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000001110001001) && ({row_reg, col_reg}<16'b1000001110001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001110001100) && ({row_reg, col_reg}<16'b1000001110010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000001110010001) && ({row_reg, col_reg}<16'b1000001110010011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000001110010011) && ({row_reg, col_reg}<16'b1000001110100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000001110100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000001110100001) && ({row_reg, col_reg}<16'b1000001110100100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001110100100) && ({row_reg, col_reg}<16'b1000001110100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000001110100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000001110100111) && ({row_reg, col_reg}<16'b1000001110101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001110101001) && ({row_reg, col_reg}<16'b1000001110111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001110111000) && ({row_reg, col_reg}<16'b1000001110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000001110111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000001110111011) && ({row_reg, col_reg}<16'b1000001110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001110111101) && ({row_reg, col_reg}<16'b1000001111000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000001111000000) && ({row_reg, col_reg}<16'b1000001111000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001111000010) && ({row_reg, col_reg}<16'b1000001111000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000001111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001111001000) && ({row_reg, col_reg}<16'b1000001111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000001111001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001111001100) && ({row_reg, col_reg}<16'b1000001111001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001111001110) && ({row_reg, col_reg}<16'b1000001111010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001111010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000001111010001) && ({row_reg, col_reg}<16'b1000001111101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000001111101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000001111110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000001111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001111110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000001111110011) && ({row_reg, col_reg}<16'b1000001111110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001111110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000001111110111) && ({row_reg, col_reg}<16'b1000001111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000001111111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000001111111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000001111111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001111111100) && ({row_reg, col_reg}<16'b1000001111111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b1000001111111110) && ({row_reg, col_reg}<16'b1000010000000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000010000000000) && ({row_reg, col_reg}<16'b1000010000000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010000000010) && ({row_reg, col_reg}<16'b1000010000001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010000001010) && ({row_reg, col_reg}<16'b1000010000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010000001100) && ({row_reg, col_reg}<16'b1000010000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000010000010010) && ({row_reg, col_reg}<16'b1000010000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000010000100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000010000100110) && ({row_reg, col_reg}<16'b1000010000101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010000101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000010000110000) && ({row_reg, col_reg}<16'b1000010000110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010000110011) && ({row_reg, col_reg}<16'b1000010000110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000010000110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000010000110110) && ({row_reg, col_reg}<16'b1000010000111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010000111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000010000111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000010000111101) && ({row_reg, col_reg}<16'b1000010000111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010000111111) && ({row_reg, col_reg}<16'b1000010001000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000010001000111) && ({row_reg, col_reg}<16'b1000010001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010001001001) && ({row_reg, col_reg}<16'b1000010001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010001010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010001010001) && ({row_reg, col_reg}<16'b1000010001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000010001010100) && ({row_reg, col_reg}<16'b1000010001011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000010001011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010001011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010001011010) && ({row_reg, col_reg}<16'b1000010001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000010001011111) && ({row_reg, col_reg}<16'b1000010001100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010001100010) && ({row_reg, col_reg}<16'b1000010001100100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010001100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000010001100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b1000010001100110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b1000010001100111) && ({row_reg, col_reg}<16'b1000010001101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000010001101001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000010001101010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010001101011) && ({row_reg, col_reg}<16'b1000010001101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000010001101111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010001110000) && ({row_reg, col_reg}<16'b1000010001110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010001110010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010001110011) && ({row_reg, col_reg}<16'b1000010001111000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000010001111000) && ({row_reg, col_reg}<16'b1000010001111011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000010001111011) && ({row_reg, col_reg}<16'b1000010010000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000010010000011) && ({row_reg, col_reg}<16'b1000010010000111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000010010000111) && ({row_reg, col_reg}<16'b1000010010001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000010010001001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000010010001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010010001011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000010010001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010010001101) && ({row_reg, col_reg}<16'b1000010010010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000010010010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000010010010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010010010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000010010010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010010010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000010010010101) && ({row_reg, col_reg}<16'b1000010010011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000010010011111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000010010100000) && ({row_reg, col_reg}<16'b1000010010100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010010100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000010010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000010010100100) && ({row_reg, col_reg}<16'b1000010010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010010101000) && ({row_reg, col_reg}<16'b1000010010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000010010110011) && ({row_reg, col_reg}<16'b1000010010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010010110101) && ({row_reg, col_reg}<16'b1000010010111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000010010111010) && ({row_reg, col_reg}<16'b1000010010111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000010010111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000010010111101) && ({row_reg, col_reg}<16'b1000010010111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010010111111) && ({row_reg, col_reg}<16'b1000010011000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000010011000001) && ({row_reg, col_reg}<16'b1000010011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010011001000) && ({row_reg, col_reg}<16'b1000010011001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000010011001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010011010000) && ({row_reg, col_reg}<16'b1000010011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000010011101110) && ({row_reg, col_reg}<16'b1000010011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000010011110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010011110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000010011110010) && ({row_reg, col_reg}<16'b1000010011110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010011110100) && ({row_reg, col_reg}<16'b1000010011111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000010011111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010011111011) && ({row_reg, col_reg}<16'b1000010011111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b1000010011111110) && ({row_reg, col_reg}<16'b1000010100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000010100010010) && ({row_reg, col_reg}<16'b1000010100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000010100100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000010100100110) && ({row_reg, col_reg}<16'b1000010100101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010100101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000010100101001) && ({row_reg, col_reg}<16'b1000010100101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000010100101011) && ({row_reg, col_reg}<16'b1000010100110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010100110001) && ({row_reg, col_reg}<16'b1000010100110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010100110111) && ({row_reg, col_reg}<16'b1000010100111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010100111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000010100111110) && ({row_reg, col_reg}<16'b1000010101000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010101000000) && ({row_reg, col_reg}<16'b1000010101010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000010101010101) && ({row_reg, col_reg}<16'b1000010101011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010101011011) && ({row_reg, col_reg}<16'b1000010101011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000010101011101) && ({row_reg, col_reg}<16'b1000010101100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010101100000) && ({row_reg, col_reg}<16'b1000010101100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010101100011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b1000010101100100) && ({row_reg, col_reg}<16'b1000010101100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000010101100110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b1000010101100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000010101101000) && ({row_reg, col_reg}<16'b1000010101101010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010101101010) && ({row_reg, col_reg}<16'b1000010101110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000010101110000) && ({row_reg, col_reg}<16'b1000010101110010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010101110010) && ({row_reg, col_reg}<16'b1000010101111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000010101111100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000010101111101) && ({row_reg, col_reg}<16'b1000010110000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000010110000010) && ({row_reg, col_reg}<16'b1000010110001010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000010110001010) && ({row_reg, col_reg}<16'b1000010110001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000010110001101) && ({row_reg, col_reg}<16'b1000010110010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000010110010000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000010110010001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000010110010010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010110010011) && ({row_reg, col_reg}<16'b1000010110011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000010110011001) && ({row_reg, col_reg}<16'b1000010110011011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b1000010110011011) && ({row_reg, col_reg}<16'b1000010110011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000010110011101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010110011110) && ({row_reg, col_reg}<16'b1000010110100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000010110100000) && ({row_reg, col_reg}<16'b1000010110100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010110100011) && ({row_reg, col_reg}<16'b1000010110101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010110101111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000010110110000) && ({row_reg, col_reg}<16'b1000010110110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000010110110010) && ({row_reg, col_reg}<16'b1000010110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010110110101) && ({row_reg, col_reg}<16'b1000010110111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010110111011) && ({row_reg, col_reg}<16'b1000010110111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000010110111101) && ({row_reg, col_reg}<16'b1000010111000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010111000110) && ({row_reg, col_reg}<16'b1000010111010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000010111010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000010111010001) && ({row_reg, col_reg}<16'b1000010111101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000010111101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000010111101110) && ({row_reg, col_reg}<16'b1000010111110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010111110001) && ({row_reg, col_reg}<16'b1000010111110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000010111110011) && ({row_reg, col_reg}<16'b1000010111110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010111110101) && ({row_reg, col_reg}<16'b1000010111110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000010111110111) && ({row_reg, col_reg}<16'b1000010111111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000010111111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010111111011) && ({row_reg, col_reg}<16'b1000010111111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b1000010111111110) && ({row_reg, col_reg}<16'b1000011000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000011000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000011000010010) && ({row_reg, col_reg}<16'b1000011000100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000011000100100) && ({row_reg, col_reg}<16'b1000011000100110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000011000100110) && ({row_reg, col_reg}<16'b1000011000101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011000101001) && ({row_reg, col_reg}<16'b1000011000101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000011000101011) && ({row_reg, col_reg}<16'b1000011000111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011000111001) && ({row_reg, col_reg}<16'b1000011000111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011000111101) && ({row_reg, col_reg}<16'b1000011001000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011001000000) && ({row_reg, col_reg}<16'b1000011001000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000011001000010) && ({row_reg, col_reg}<16'b1000011001010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000011001010111) && ({row_reg, col_reg}<16'b1000011001011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000011001011011) && ({row_reg, col_reg}<16'b1000011001011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000011001011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000011001011110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1000011001011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000011001100000) && ({row_reg, col_reg}<16'b1000011001100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000011001100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b1000011001100100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b1000011001100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b1000011001100110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b1000011001100111) && ({row_reg, col_reg}<16'b1000011001110100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000011001110100) && ({row_reg, col_reg}<16'b1000011001110110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b1000011001110110) && ({row_reg, col_reg}<16'b1000011001111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000011001111101) && ({row_reg, col_reg}<16'b1000011001111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000011001111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000011010000000) && ({row_reg, col_reg}<16'b1000011010000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000011010000011) && ({row_reg, col_reg}<16'b1000011010000101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b1000011010000101) && ({row_reg, col_reg}<16'b1000011010001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000011010001011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000011010001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000011010001101) && ({row_reg, col_reg}<16'b1000011010011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000011010011100) && ({row_reg, col_reg}<16'b1000011010011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000011010011110) && ({row_reg, col_reg}<16'b1000011010100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000011010100011) && ({row_reg, col_reg}<16'b1000011010101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000011010101100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000011010101101) && ({row_reg, col_reg}<16'b1000011010101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000011010101111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000011010110000) && ({row_reg, col_reg}<16'b1000011010111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000011010111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000011010111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011010111011) && ({row_reg, col_reg}<16'b1000011010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011010111110) && ({row_reg, col_reg}<16'b1000011011010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000011011010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000011011010001) && ({row_reg, col_reg}<16'b1000011011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000011011101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000011011101110) && ({row_reg, col_reg}<16'b1000011011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000011011110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011011110001) && ({row_reg, col_reg}<16'b1000011011110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000011011110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000011011110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000011011110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000011011110110) && ({row_reg, col_reg}<16'b1000011011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011011111011) && ({row_reg, col_reg}<16'b1000011011111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b1000011011111110) && ({row_reg, col_reg}<16'b1000011100001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011100001001) && ({row_reg, col_reg}<16'b1000011100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011100001011) && ({row_reg, col_reg}<16'b1000011100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000011100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000011100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011100010010) && ({row_reg, col_reg}<16'b1000011100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000011100100011) && ({row_reg, col_reg}<16'b1000011100100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000011100100101) && ({row_reg, col_reg}<16'b1000011100101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011100101001) && ({row_reg, col_reg}<16'b1000011100101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000011100101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000011100101101) && ({row_reg, col_reg}<16'b1000011100101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000011100101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000011100110000) && ({row_reg, col_reg}<16'b1000011100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000011100110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000011100110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000011100110101) && ({row_reg, col_reg}<16'b1000011100111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000011100111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000011100111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000011100111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011100111100) && ({row_reg, col_reg}<16'b1000011101000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011101000010) && ({row_reg, col_reg}<16'b1000011101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000011101000100) && ({row_reg, col_reg}<16'b1000011101000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000011101000111) && ({row_reg, col_reg}<16'b1000011101001001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000011101001001) && ({row_reg, col_reg}<16'b1000011101011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000011101011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000011101011110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000011101011111) && ({row_reg, col_reg}<16'b1000011101100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000011101100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b1000011101100100) && ({row_reg, col_reg}<16'b1000011101100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b1000011101100111) && ({row_reg, col_reg}<16'b1000011101111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000011101111101) && ({row_reg, col_reg}<16'b1000011101111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000011101111111) && ({row_reg, col_reg}<16'b1000011110000010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000011110000010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b1000011110000011) && ({row_reg, col_reg}<16'b1000011110000101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b1000011110000101) && ({row_reg, col_reg}<16'b1000011110011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000011110011001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000011110011010) && ({row_reg, col_reg}<16'b1000011110011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000011110011101) && ({row_reg, col_reg}<16'b1000011110100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000011110100010) && ({row_reg, col_reg}<16'b1000011110100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000011110100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000011110100111) && ({row_reg, col_reg}<16'b1000011110101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000011110101011) && ({row_reg, col_reg}<16'b1000011110101101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000011110101101) && ({row_reg, col_reg}<16'b1000011110110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000011110110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000011110111000) && ({row_reg, col_reg}<16'b1000011110111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011110111010) && ({row_reg, col_reg}<16'b1000011110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011110111101) && ({row_reg, col_reg}<16'b1000011111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011111000000) && ({row_reg, col_reg}<16'b1000011111000010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000011111000010) && ({row_reg, col_reg}<16'b1000011111001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011111001010) && ({row_reg, col_reg}<16'b1000011111001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000011111001100) && ({row_reg, col_reg}<16'b1000011111001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011111001110) && ({row_reg, col_reg}<16'b1000011111010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011111010000) && ({row_reg, col_reg}<16'b1000011111010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000011111010010) && ({row_reg, col_reg}<16'b1000011111101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000011111101110) && ({row_reg, col_reg}<16'b1000011111110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011111110000) && ({row_reg, col_reg}<16'b1000011111110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000011111110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000011111110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000011111110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000011111110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011111110111) && ({row_reg, col_reg}<16'b1000011111111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011111111011) && ({row_reg, col_reg}<16'b1000011111111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000011111111110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}==16'b1000011111111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100000000000) && ({row_reg, col_reg}<16'b1000100000001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100000001000) && ({row_reg, col_reg}<16'b1000100000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100000001100) && ({row_reg, col_reg}<16'b1000100000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100000010000) && ({row_reg, col_reg}<16'b1000100000010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000100000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100000010011) && ({row_reg, col_reg}<16'b1000100000010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100000010101) && ({row_reg, col_reg}<16'b1000100000011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100000011001) && ({row_reg, col_reg}<16'b1000100000011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100000011101) && ({row_reg, col_reg}<16'b1000100000011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100000011111) && ({row_reg, col_reg}<16'b1000100000100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100000100011) && ({row_reg, col_reg}<16'b1000100000101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100000101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100000101010) && ({row_reg, col_reg}<16'b1000100000101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000100000101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000100000101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1000100000101111)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b1000100000110000) && ({row_reg, col_reg}<16'b1000100000110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000100000110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000100000110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000100000110101) && ({row_reg, col_reg}<16'b1000100000111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100000111000) && ({row_reg, col_reg}<16'b1000100000111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000100000111010) && ({row_reg, col_reg}<16'b1000100000111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000100000111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000100000111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000100000111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000100000111111) && ({row_reg, col_reg}<16'b1000100001000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100001000001) && ({row_reg, col_reg}<16'b1000100001000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000100001000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000100001000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000100001000110) && ({row_reg, col_reg}<16'b1000100001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000100001011111) && ({row_reg, col_reg}<16'b1000100001100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000100001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100001100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000100001100100) && ({row_reg, col_reg}<16'b1000100001100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b1000100001100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000100001101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b1000100001101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100001101010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000100001101011) && ({row_reg, col_reg}<16'b1000100001111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000100001111101) && ({row_reg, col_reg}<16'b1000100001111111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000100001111111) && ({row_reg, col_reg}<16'b1000100010000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000100010000011) && ({row_reg, col_reg}<16'b1000100010000110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b1000100010000110) && ({row_reg, col_reg}<16'b1000100010010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000100010010100) && ({row_reg, col_reg}<16'b1000100010010110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000100010010110) && ({row_reg, col_reg}<16'b1000100010011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100010011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000100010011010) && ({row_reg, col_reg}<16'b1000100010011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000100010011100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000100010011101) && ({row_reg, col_reg}<16'b1000100010011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000100010011111) && ({row_reg, col_reg}<16'b1000100010110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100010110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000100010110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000100010111000) && ({row_reg, col_reg}<16'b1000100010111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100010111100) && ({row_reg, col_reg}<16'b1000100010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000100010111111)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b1000100011000000) && ({row_reg, col_reg}<16'b1000100011000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000100011000010) && ({row_reg, col_reg}<16'b1000100011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000100011001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1000100011001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000100011001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100011001101) && ({row_reg, col_reg}<16'b1000100011010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100011010010) && ({row_reg, col_reg}<16'b1000100011010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100011010100) && ({row_reg, col_reg}<16'b1000100011011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100011011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100011011010) && ({row_reg, col_reg}<16'b1000100011011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100011011100) && ({row_reg, col_reg}<16'b1000100011100100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100011100100) && ({row_reg, col_reg}<16'b1000100011101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100011101001) && ({row_reg, col_reg}<16'b1000100011101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100011101011) && ({row_reg, col_reg}<16'b1000100011110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000100011110011) && ({row_reg, col_reg}<16'b1000100011110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100011110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100011110110) && ({row_reg, col_reg}<16'b1000100011111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000100011111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100011111011) && ({row_reg, col_reg}<16'b1000100011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000100011111110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}==16'b1000100011111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000100100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100100000001) && ({row_reg, col_reg}<16'b1000100100001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100100001001) && ({row_reg, col_reg}<16'b1000100100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100100001011) && ({row_reg, col_reg}<16'b1000100100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100100010001) && ({row_reg, col_reg}<16'b1000100100010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100100010011) && ({row_reg, col_reg}<16'b1000100100101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100100101000) && ({row_reg, col_reg}<16'b1000100100101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000100100101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100100101100) && ({row_reg, col_reg}<16'b1000100100110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000100100110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000100100111000) && ({row_reg, col_reg}<16'b1000100100111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000100100111010) && ({row_reg, col_reg}<16'b1000100100111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100100111100) && ({row_reg, col_reg}<16'b1000100100111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000100100111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000100100111111) && ({row_reg, col_reg}<16'b1000100101000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000100101000010) && ({row_reg, col_reg}<16'b1000100101000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100101000100) && ({row_reg, col_reg}<16'b1000100101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000100101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000100101000111) && ({row_reg, col_reg}<16'b1000100101010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000100101010001) && ({row_reg, col_reg}<16'b1000100101010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000100101010011) && ({row_reg, col_reg}<16'b1000100101100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100101100000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b1000100101100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1000100101100010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b1000100101100011)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b1000100101100100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b1000100101100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b1000100101100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000100101100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b1000100101101000) && ({row_reg, col_reg}<16'b1000100101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000100101101010) && ({row_reg, col_reg}<16'b1000100101101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100101101100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000100101101101) && ({row_reg, col_reg}<16'b1000100110010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000100110010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000100110010101) && ({row_reg, col_reg}<16'b1000100110010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100110010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000100110011000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000100110011001) && ({row_reg, col_reg}<16'b1000100110011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000100110011100) && ({row_reg, col_reg}<16'b1000100110011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000100110011111) && ({row_reg, col_reg}<16'b1000100110110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100110110001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000100110110010) && ({row_reg, col_reg}<16'b1000100110110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000100110110110) && ({row_reg, col_reg}<16'b1000100110111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000100110111000) && ({row_reg, col_reg}<16'b1000100110111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100110111010) && ({row_reg, col_reg}<16'b1000100110111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000100110111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000100110111101) && ({row_reg, col_reg}<16'b1000100110111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100110111111) && ({row_reg, col_reg}<16'b1000100111000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1000100111000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000100111000101) && ({row_reg, col_reg}<16'b1000100111000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100111000111) && ({row_reg, col_reg}<16'b1000100111001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000100111001001) && ({row_reg, col_reg}<16'b1000100111001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100111001100) && ({row_reg, col_reg}<16'b1000100111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100111010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100111010010) && ({row_reg, col_reg}<16'b1000100111100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100111100100) && ({row_reg, col_reg}<16'b1000100111100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100111100110) && ({row_reg, col_reg}<16'b1000100111101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100111101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100111101010) && ({row_reg, col_reg}<16'b1000100111110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000100111110011) && ({row_reg, col_reg}<16'b1000100111110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100111110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100111110110) && ({row_reg, col_reg}<16'b1000100111111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100111111001) && ({row_reg, col_reg}<16'b1000100111111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100111111011) && ({row_reg, col_reg}<16'b1000100111111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000100111111110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}==16'b1000100111111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101000000000) && ({row_reg, col_reg}<16'b1000101000001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101000001010) && ({row_reg, col_reg}<16'b1000101000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101000001100) && ({row_reg, col_reg}<16'b1000101000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000101000001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101000010000) && ({row_reg, col_reg}<16'b1000101000100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101000100101) && ({row_reg, col_reg}<16'b1000101000101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000101000101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101000101001) && ({row_reg, col_reg}<16'b1000101000101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101000101100) && ({row_reg, col_reg}<16'b1000101000101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101000101110) && ({row_reg, col_reg}<16'b1000101000110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101000110110) && ({row_reg, col_reg}<16'b1000101000111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000101000111001) && ({row_reg, col_reg}<16'b1000101000111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101000111100) && ({row_reg, col_reg}<16'b1000101000111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1000101000111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000101000111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000101001000000) && ({row_reg, col_reg}<16'b1000101001000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101001000010) && ({row_reg, col_reg}<16'b1000101001000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101001000101) && ({row_reg, col_reg}<16'b1000101001001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000101001001000) && ({row_reg, col_reg}<16'b1000101001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101001001011) && ({row_reg, col_reg}<16'b1000101001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000101001010000) && ({row_reg, col_reg}<16'b1000101001010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000101001010100) && ({row_reg, col_reg}<16'b1000101001011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000101001011110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b1000101001011111) && ({row_reg, col_reg}<16'b1000101001100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b1000101001100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000101001100100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b1000101001100101) && ({row_reg, col_reg}<16'b1000101001100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000101001100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000101001101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000101001101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000101001101010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1000101001101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101001101100) && ({row_reg, col_reg}<16'b1000101001110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000101001110000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000101001110001) && ({row_reg, col_reg}<16'b1000101010001010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000101010001010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b1000101010001011) && ({row_reg, col_reg}<16'b1000101010010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000101010010010) && ({row_reg, col_reg}<16'b1000101010010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000101010010110) && ({row_reg, col_reg}<16'b1000101010011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101010011000) && ({row_reg, col_reg}<16'b1000101010011011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000101010011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101010011100) && ({row_reg, col_reg}<16'b1000101010110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000101010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101010110101) && ({row_reg, col_reg}<16'b1000101010111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000101010111001) && ({row_reg, col_reg}<16'b1000101010111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101010111011) && ({row_reg, col_reg}<16'b1000101010111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000101010111101) && ({row_reg, col_reg}<16'b1000101010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000101010111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101011000000) && ({row_reg, col_reg}<16'b1000101011000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1000101011000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000101011000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000101011000101)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==16'b1000101011000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000101011000111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000101011001000) && ({row_reg, col_reg}<16'b1000101011001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000101011001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101011001101) && ({row_reg, col_reg}<16'b1000101011001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000101011001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101011010000) && ({row_reg, col_reg}<16'b1000101011010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101011010010) && ({row_reg, col_reg}<16'b1000101011100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101011100000) && ({row_reg, col_reg}<16'b1000101011100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101011100010) && ({row_reg, col_reg}<16'b1000101011101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000101011101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101011101011) && ({row_reg, col_reg}<16'b1000101011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000101011110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101011110011) && ({row_reg, col_reg}<16'b1000101011110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000101011110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101011110110) && ({row_reg, col_reg}<16'b1000101011111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000101011111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101011111010) && ({row_reg, col_reg}<16'b1000101011111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101011111100) && ({row_reg, col_reg}<16'b1000101011111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000101011111110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}==16'b1000101011111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101100000000) && ({row_reg, col_reg}<16'b1000101100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101100000101) && ({row_reg, col_reg}<16'b1000101100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101100000111) && ({row_reg, col_reg}<16'b1000101100001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000101100001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101100001010) && ({row_reg, col_reg}<16'b1000101100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101100001100) && ({row_reg, col_reg}<16'b1000101100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000101100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101100010000) && ({row_reg, col_reg}<16'b1000101100100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101100100101) && ({row_reg, col_reg}<16'b1000101100101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101100101000) && ({row_reg, col_reg}<16'b1000101100101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000101100101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101100101101) && ({row_reg, col_reg}<16'b1000101100101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101100101111) && ({row_reg, col_reg}<16'b1000101100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101100110110) && ({row_reg, col_reg}<16'b1000101100111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000101100111001) && ({row_reg, col_reg}<16'b1000101100111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000101100111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000101100111101) && ({row_reg, col_reg}<16'b1000101100111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000101100111111) && ({row_reg, col_reg}<16'b1000101101000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000101101000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101101000011) && ({row_reg, col_reg}<16'b1000101101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000101101000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101101000111) && ({row_reg, col_reg}<16'b1000101101001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000101101001100) && ({row_reg, col_reg}<16'b1000101101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000101101010000) && ({row_reg, col_reg}<16'b1000101101010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000101101010011) && ({row_reg, col_reg}<16'b1000101101011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000101101011001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000101101011010) && ({row_reg, col_reg}<16'b1000101101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000101101011110) && ({row_reg, col_reg}<16'b1000101101100010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b1000101101100010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b1000101101100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000101101100100) && ({row_reg, col_reg}<16'b1000101101100110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000101101100110) && ({row_reg, col_reg}<16'b1000101101101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000101101101000) && ({row_reg, col_reg}<16'b1000101101110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000101101110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000101101110001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000101101110010) && ({row_reg, col_reg}<16'b1000101110010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000101110010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000101110010001) && ({row_reg, col_reg}<16'b1000101110010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000101110010011) && ({row_reg, col_reg}<16'b1000101110011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101110011010) && ({row_reg, col_reg}<16'b1000101110100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000101110100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000101110100001) && ({row_reg, col_reg}<16'b1000101110110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000101110110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000101110110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000101110110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101110110101) && ({row_reg, col_reg}<16'b1000101110111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000101110111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000101110111001) && ({row_reg, col_reg}<16'b1000101110111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101110111011) && ({row_reg, col_reg}<16'b1000101110111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000101110111101) && ({row_reg, col_reg}<16'b1000101111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000101111000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000101111000001) && ({row_reg, col_reg}<16'b1000101111000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000101111000011) && ({row_reg, col_reg}<16'b1000101111000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101111000101) && ({row_reg, col_reg}<16'b1000101111000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101111000111) && ({row_reg, col_reg}<16'b1000101111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000101111001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101111001100) && ({row_reg, col_reg}<16'b1000101111001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101111001110) && ({row_reg, col_reg}<16'b1000101111010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101111010000) && ({row_reg, col_reg}<16'b1000101111010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101111010011) && ({row_reg, col_reg}<16'b1000101111100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101111100000) && ({row_reg, col_reg}<16'b1000101111100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101111100011) && ({row_reg, col_reg}<16'b1000101111101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000101111101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101111101011) && ({row_reg, col_reg}<16'b1000101111101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000101111101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000101111101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101111101111) && ({row_reg, col_reg}<16'b1000101111110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000101111110010) && ({row_reg, col_reg}<16'b1000101111110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101111110100) && ({row_reg, col_reg}<16'b1000101111111111)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}==16'b1000101111111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000110000000000) && ({row_reg, col_reg}<16'b1000110000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110000000110) && ({row_reg, col_reg}<16'b1000110000001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110000001000) && ({row_reg, col_reg}<16'b1000110000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110000001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000110000010000) && ({row_reg, col_reg}<16'b1000110000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110000010010) && ({row_reg, col_reg}<16'b1000110000011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110000011001) && ({row_reg, col_reg}<16'b1000110000011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110000011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000110000011100) && ({row_reg, col_reg}<16'b1000110000101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110000101101) && ({row_reg, col_reg}<16'b1000110000101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000110000101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110000110000) && ({row_reg, col_reg}<16'b1000110000110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110000110011) && ({row_reg, col_reg}<16'b1000110000111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000110000111100) && ({row_reg, col_reg}<16'b1000110001000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110001000010) && ({row_reg, col_reg}<16'b1000110001001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110001001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000110001001001) && ({row_reg, col_reg}<16'b1000110001001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110001001100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000110001001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110001001110) && ({row_reg, col_reg}<16'b1000110001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110001010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110001010001) && ({row_reg, col_reg}<16'b1000110001010011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000110001010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110001010100) && ({row_reg, col_reg}<16'b1000110001011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000110001011000) && ({row_reg, col_reg}<16'b1000110001011010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110001011010) && ({row_reg, col_reg}<16'b1000110001011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110001011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000110001011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000110001011111) && ({row_reg, col_reg}<16'b1000110001100010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b1000110001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110001100011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000110001100100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000110001100101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110001100110) && ({row_reg, col_reg}<16'b1000110001101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110001101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000110001101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000110001101011) && ({row_reg, col_reg}<16'b1000110001101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110001101101) && ({row_reg, col_reg}<16'b1000110001101111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1000110001101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000110001110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110001110001) && ({row_reg, col_reg}<16'b1000110001110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000110001110101) && ({row_reg, col_reg}<16'b1000110001111000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000110001111000) && ({row_reg, col_reg}<16'b1000110001111010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b1000110001111010) && ({row_reg, col_reg}<16'b1000110001111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000110001111101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000110001111110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110001111111) && ({row_reg, col_reg}<16'b1000110010000011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000110010000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000110010000100) && ({row_reg, col_reg}<16'b1000110010000111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110010000111) && ({row_reg, col_reg}<16'b1000110010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000110010001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000110010001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110010001110) && ({row_reg, col_reg}<16'b1000110010010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110010010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110010010010) && ({row_reg, col_reg}<16'b1000110010010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000110010010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110010010101) && ({row_reg, col_reg}<16'b1000110010010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000110010010111) && ({row_reg, col_reg}<16'b1000110010011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110010011001) && ({row_reg, col_reg}<16'b1000110010011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110010011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000110010011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000110010011111) && ({row_reg, col_reg}<16'b1000110010100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110010100001) && ({row_reg, col_reg}<16'b1000110010101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000110010101001) && ({row_reg, col_reg}<16'b1000110010101100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110010101100) && ({row_reg, col_reg}<16'b1000110010110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110010110001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000110010110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000110010110011) && ({row_reg, col_reg}<16'b1000110010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110010110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000110010110111) && ({row_reg, col_reg}<16'b1000110010111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000110010111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000110010111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000110010111011) && ({row_reg, col_reg}<16'b1000110010111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110010111101) && ({row_reg, col_reg}<16'b1000110010111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000110010111111) && ({row_reg, col_reg}<16'b1000110011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000110011000001)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==16'b1000110011000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000110011000011) && ({row_reg, col_reg}<16'b1000110011000101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000110011000101) && ({row_reg, col_reg}<16'b1000110011000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000110011000111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000110011001000) && ({row_reg, col_reg}<16'b1000110011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000110011001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110011001100) && ({row_reg, col_reg}<16'b1000110011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000110011001110) && ({row_reg, col_reg}<16'b1000110011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110011010001) && ({row_reg, col_reg}<16'b1000110011010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110011010111) && ({row_reg, col_reg}<16'b1000110011101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110011101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110011101100) && ({row_reg, col_reg}<16'b1000110011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110011101111) && ({row_reg, col_reg}<16'b1000110011110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110011110001) && ({row_reg, col_reg}<16'b1000110011110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110011110111)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b1000110011111000) && ({row_reg, col_reg}<16'b1000110100000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110100000111) && ({row_reg, col_reg}<16'b1000110100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110100001001) && ({row_reg, col_reg}<16'b1000110100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000110100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110100010001) && ({row_reg, col_reg}<16'b1000110100011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110100011001) && ({row_reg, col_reg}<16'b1000110100101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110100101110) && ({row_reg, col_reg}<16'b1000110100110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000110100110000) && ({row_reg, col_reg}<16'b1000110100110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110100110011) && ({row_reg, col_reg}<16'b1000110100110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000110100110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000110100110110) && ({row_reg, col_reg}<16'b1000110100111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000110100111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110100111101) && ({row_reg, col_reg}<16'b1000110100111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110100111111) && ({row_reg, col_reg}<16'b1000110101000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000110101000001) && ({row_reg, col_reg}<16'b1000110101001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000110101001001) && ({row_reg, col_reg}<16'b1000110101001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110101001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000110101001110) && ({row_reg, col_reg}<16'b1000110101010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110101010000) && ({row_reg, col_reg}<16'b1000110101011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000110101011000) && ({row_reg, col_reg}<16'b1000110101011010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110101011010) && ({row_reg, col_reg}<16'b1000110101100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110101100000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b1000110101100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110101100010) && ({row_reg, col_reg}<16'b1000110101100100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110101100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000110101100101) && ({row_reg, col_reg}<16'b1000110101101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000110101101100) && ({row_reg, col_reg}<16'b1000110101101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000110101101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000110101110000) && ({row_reg, col_reg}<16'b1000110101110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000110101110010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000110101110011) && ({row_reg, col_reg}<16'b1000110101110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110101110101) && ({row_reg, col_reg}<16'b1000110101111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000110101111000) && ({row_reg, col_reg}<16'b1000110101111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000110101111101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000110101111110) && ({row_reg, col_reg}<16'b1000110110000001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110110000001) && ({row_reg, col_reg}<16'b1000110110000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000110110000100) && ({row_reg, col_reg}<16'b1000110110000111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110110000111) && ({row_reg, col_reg}<16'b1000110110001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000110110001001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110110001010) && ({row_reg, col_reg}<16'b1000110110001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000110110001111) && ({row_reg, col_reg}<16'b1000110110010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110110010001) && ({row_reg, col_reg}<16'b1000110110010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000110110010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110110010101) && ({row_reg, col_reg}<16'b1000110110011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000110110011100) && ({row_reg, col_reg}<16'b1000110110100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110110100001) && ({row_reg, col_reg}<16'b1000110110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000110110100111) && ({row_reg, col_reg}<16'b1000110110101001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110110101001) && ({row_reg, col_reg}<16'b1000110110110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000110110110000) && ({row_reg, col_reg}<16'b1000110110110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000110110110010) && ({row_reg, col_reg}<16'b1000110110110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110110110101) && ({row_reg, col_reg}<16'b1000110110110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000110110110111) && ({row_reg, col_reg}<16'b1000110110111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000110110111010) && ({row_reg, col_reg}<16'b1000110110111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000110110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000110111000000) && ({row_reg, col_reg}<16'b1000110111000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000110111000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000110111000011) && ({row_reg, col_reg}<16'b1000110111000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000110111000101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000110111000110) && ({row_reg, col_reg}<16'b1000110111001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000110111001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000110111001001) && ({row_reg, col_reg}<16'b1000110111001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110111001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000110111001100) && ({row_reg, col_reg}<16'b1000110111010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110111010010) && ({row_reg, col_reg}<16'b1000110111011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110111011000) && ({row_reg, col_reg}<16'b1000110111100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110111100000) && ({row_reg, col_reg}<16'b1000110111100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110111100010) && ({row_reg, col_reg}<16'b1000110111101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110111101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110111101100) && ({row_reg, col_reg}<16'b1000110111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110111101111) && ({row_reg, col_reg}<16'b1000110111111000)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b1000110111111000) && ({row_reg, col_reg}<16'b1000111000001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111000001000) && ({row_reg, col_reg}<16'b1000111000001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111000001010) && ({row_reg, col_reg}<16'b1000111000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111000010001) && ({row_reg, col_reg}<16'b1000111000010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111000010011) && ({row_reg, col_reg}<16'b1000111000011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111000011000) && ({row_reg, col_reg}<16'b1000111000011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111000011011) && ({row_reg, col_reg}<16'b1000111000101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000111000101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000111000110000) && ({row_reg, col_reg}<16'b1000111000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000111000110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000111000110101) && ({row_reg, col_reg}<16'b1000111000111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111000111001) && ({row_reg, col_reg}<16'b1000111000111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000111000111011) && ({row_reg, col_reg}<16'b1000111000111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000111000111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111000111110) && ({row_reg, col_reg}<16'b1000111001000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000111001000000) && ({row_reg, col_reg}<16'b1000111001000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111001000100) && ({row_reg, col_reg}<16'b1000111001000111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000111001000111) && ({row_reg, col_reg}<16'b1000111001001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000111001001010) && ({row_reg, col_reg}<16'b1000111001001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111001001110) && ({row_reg, col_reg}<16'b1000111001010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000111001010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111001010001) && ({row_reg, col_reg}<16'b1000111001011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111001011000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000111001011001) && ({row_reg, col_reg}<16'b1000111001100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111001100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000111001100100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b1000111001100101) && ({row_reg, col_reg}<16'b1000111001101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111001101000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000111001101001) && ({row_reg, col_reg}<16'b1000111001101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000111001101100) && ({row_reg, col_reg}<16'b1000111001101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111001101110) && ({row_reg, col_reg}<16'b1000111001110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000111001110000) && ({row_reg, col_reg}<16'b1000111001110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111001110101) && ({row_reg, col_reg}<16'b1000111001110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000111001110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111001111000) && ({row_reg, col_reg}<16'b1000111001111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000111001111011) && ({row_reg, col_reg}<16'b1000111001111101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000111001111101) && ({row_reg, col_reg}<16'b1000111001111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000111001111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000111010000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111010000001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000111010000010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000111010000011) && ({row_reg, col_reg}<16'b1000111010001000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000111010001000) && ({row_reg, col_reg}<16'b1000111010001010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000111010001010) && ({row_reg, col_reg}<16'b1000111010001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000111010001100) && ({row_reg, col_reg}<16'b1000111010010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111010010011) && ({row_reg, col_reg}<16'b1000111010010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000111010010110) && ({row_reg, col_reg}<16'b1000111010011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111010011000) && ({row_reg, col_reg}<16'b1000111010011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000111010011100) && ({row_reg, col_reg}<16'b1000111010100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000111010100010) && ({row_reg, col_reg}<16'b1000111010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111010100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000111010101000) && ({row_reg, col_reg}<16'b1000111010101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111010101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111010110000) && ({row_reg, col_reg}<16'b1000111010110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000111010110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111010110011) && ({row_reg, col_reg}<16'b1000111010110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000111010110111) && ({row_reg, col_reg}<16'b1000111010111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000111010111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111010111010) && ({row_reg, col_reg}<16'b1000111010111100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000111010111100) && ({row_reg, col_reg}<16'b1000111011000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111011000000) && ({row_reg, col_reg}<16'b1000111011000010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000111011000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1000111011000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111011000100) && ({row_reg, col_reg}<16'b1000111011000110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000111011000110) && ({row_reg, col_reg}<16'b1000111011001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000111011001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111011001001) && ({row_reg, col_reg}<16'b1000111011001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111011001111) && ({row_reg, col_reg}<16'b1000111011010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111011010001) && ({row_reg, col_reg}<16'b1000111011011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000111011011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000111011011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111011011111) && ({row_reg, col_reg}<16'b1000111011100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111011100101) && ({row_reg, col_reg}<16'b1000111011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000111011110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111011110011) && ({row_reg, col_reg}<16'b1000111011111111)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}==16'b1000111011111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000111100000000) && ({row_reg, col_reg}<16'b1000111100001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111100001000) && ({row_reg, col_reg}<16'b1000111100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111100001010) && ({row_reg, col_reg}<16'b1000111100011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000111100011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111100011011) && ({row_reg, col_reg}<16'b1000111100101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000111100101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000111100101010) && ({row_reg, col_reg}<16'b1000111100101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111100101111) && ({row_reg, col_reg}<16'b1000111100110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000111100110010) && ({row_reg, col_reg}<16'b1000111100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000111100110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000111100110110) && ({row_reg, col_reg}<16'b1000111100111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000111100111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000111100111010) && ({row_reg, col_reg}<16'b1000111100111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111100111101) && ({row_reg, col_reg}<16'b1000111101000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000111101000000) && ({row_reg, col_reg}<16'b1000111101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111101001001) && ({row_reg, col_reg}<16'b1000111101001100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000111101001100) && ({row_reg, col_reg}<16'b1000111101010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000111101010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000111101010101) && ({row_reg, col_reg}<16'b1000111101010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111101010111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000111101011000) && ({row_reg, col_reg}<16'b1000111101100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111101100001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1000111101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111101100011) && ({row_reg, col_reg}<16'b1000111101100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000111101100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000111101100110) && ({row_reg, col_reg}<16'b1000111101101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111101101000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000111101101001) && ({row_reg, col_reg}<16'b1000111101101011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000111101101011) && ({row_reg, col_reg}<16'b1000111101110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000111101110001) && ({row_reg, col_reg}<16'b1000111101110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111101110101) && ({row_reg, col_reg}<16'b1000111101111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000111101111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111101111010) && ({row_reg, col_reg}<16'b1000111101111110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111101111110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000111101111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000111110000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111110000001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000111110000010) && ({row_reg, col_reg}<16'b1000111110000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000111110000111) && ({row_reg, col_reg}<16'b1000111110001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000111110001010) && ({row_reg, col_reg}<16'b1000111110001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000111110001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000111110001101) && ({row_reg, col_reg}<16'b1000111110001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111110001111) && ({row_reg, col_reg}<16'b1000111110101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000111110101100) && ({row_reg, col_reg}<16'b1000111110101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111110101110) && ({row_reg, col_reg}<16'b1000111110110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000111110110000) && ({row_reg, col_reg}<16'b1000111110110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000111110110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000111110110100) && ({row_reg, col_reg}<16'b1000111110110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000111110110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000111110111000) && ({row_reg, col_reg}<16'b1000111110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111110111101) && ({row_reg, col_reg}<16'b1000111110111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000111110111111) && ({row_reg, col_reg}<16'b1000111111000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000111111000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000111111000011) && ({row_reg, col_reg}<16'b1000111111000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000111111000111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000111111001000) && ({row_reg, col_reg}<16'b1000111111011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000111111011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000111111011100) && ({row_reg, col_reg}<16'b1000111111111111)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}==16'b1000111111111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001000000000000) && ({row_reg, col_reg}<16'b1001000000001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000000001000) && ({row_reg, col_reg}<16'b1001000000001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000000001010) && ({row_reg, col_reg}<16'b1001000000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000000001101) && ({row_reg, col_reg}<16'b1001000000001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001000000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000000010000) && ({row_reg, col_reg}<16'b1001000000010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001000000010011) && ({row_reg, col_reg}<16'b1001000000010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000000010110) && ({row_reg, col_reg}<16'b1001000000011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000000011000) && ({row_reg, col_reg}<16'b1001000000011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000000011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000000011101) && ({row_reg, col_reg}<16'b1001000000100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000000100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000000100010) && ({row_reg, col_reg}<16'b1001000000100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000000100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000000100111) && ({row_reg, col_reg}<16'b1001000000110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000000110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001000000110111) && ({row_reg, col_reg}<16'b1001000000111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000000111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001000000111010) && ({row_reg, col_reg}<16'b1001000001000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001000001000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000001000010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001000001000011) && ({row_reg, col_reg}<16'b1001000001000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000001000111) && ({row_reg, col_reg}<16'b1001000001001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001000001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000001001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001000001001011) && ({row_reg, col_reg}<16'b1001000001001110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001000001001110) && ({row_reg, col_reg}<16'b1001000001010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001000001010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000001010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001000001010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000001010011) && ({row_reg, col_reg}<16'b1001000001010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001000001010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000001010110) && ({row_reg, col_reg}<16'b1001000001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001000001011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000001100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001000001100001) && ({row_reg, col_reg}<16'b1001000001100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000001100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000001100100) && ({row_reg, col_reg}<16'b1001000001100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001000001100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000001100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001000001101000) && ({row_reg, col_reg}<16'b1001000001101011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001000001101011) && ({row_reg, col_reg}<16'b1001000001110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001000001110101) && ({row_reg, col_reg}<16'b1001000001111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000001111010) && ({row_reg, col_reg}<16'b1001000010000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001000010000001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001000010000010) && ({row_reg, col_reg}<16'b1001000010000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001000010000101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001000010000110) && ({row_reg, col_reg}<16'b1001000010001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001000010001000) && ({row_reg, col_reg}<16'b1001000010001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000010001010) && ({row_reg, col_reg}<16'b1001000010001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001000010001100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001000010001101) && ({row_reg, col_reg}<16'b1001000010010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001000010010010) && ({row_reg, col_reg}<16'b1001000010010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001000010010100) && ({row_reg, col_reg}<16'b1001000010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001000010100011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001000010100100) && ({row_reg, col_reg}<16'b1001000010101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001000010101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000010101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001000010101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000010101111) && ({row_reg, col_reg}<16'b1001000010110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001000010110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001000010110011) && ({row_reg, col_reg}<16'b1001000010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000010110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001000010110110) && ({row_reg, col_reg}<16'b1001000010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000010111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001000010111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000010111010) && ({row_reg, col_reg}<16'b1001000011000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001000011000000) && ({row_reg, col_reg}<16'b1001000011000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000011000010) && ({row_reg, col_reg}<16'b1001000011000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001000011000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001000011000111) && ({row_reg, col_reg}<16'b1001000011001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000011001100) && ({row_reg, col_reg}<16'b1001000011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000011110001)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b1001000011110010) && ({row_reg, col_reg}<16'b1001000100001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000100001000) && ({row_reg, col_reg}<16'b1001000100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000100001010) && ({row_reg, col_reg}<16'b1001000100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001000100010000) && ({row_reg, col_reg}<16'b1001000100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001000100010011) && ({row_reg, col_reg}<16'b1001000100010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000100010110) && ({row_reg, col_reg}<16'b1001000100011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000100011000) && ({row_reg, col_reg}<16'b1001000100011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000100011011) && ({row_reg, col_reg}<16'b1001000100011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000100011101) && ({row_reg, col_reg}<16'b1001000100100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000100100000) && ({row_reg, col_reg}<16'b1001000100100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000100100010) && ({row_reg, col_reg}<16'b1001000100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000100110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001000100110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000100110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001000100111000) && ({row_reg, col_reg}<16'b1001000100111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000100111100) && ({row_reg, col_reg}<16'b1001000100111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001000100111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000100111111)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b1001000101000000) && ({row_reg, col_reg}<16'b1001000101000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000101000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001000101000011) && ({row_reg, col_reg}<16'b1001000101000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000101000111) && ({row_reg, col_reg}<16'b1001000101001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001000101001001) && ({row_reg, col_reg}<16'b1001000101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000101001011) && ({row_reg, col_reg}<16'b1001000101001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001000101001101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001000101001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001000101001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000101010000) && ({row_reg, col_reg}<16'b1001000101010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001000101010010) && ({row_reg, col_reg}<16'b1001000101010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000101010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001000101010110) && ({row_reg, col_reg}<16'b1001000101011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000101011010) && ({row_reg, col_reg}<16'b1001000101100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001000101100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000101100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001000101100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000101100110) && ({row_reg, col_reg}<16'b1001000101101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001000101101001) && ({row_reg, col_reg}<16'b1001000101101101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001000101101101) && ({row_reg, col_reg}<16'b1001000101110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001000101110101) && ({row_reg, col_reg}<16'b1001000101110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000101110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001000101111000) && ({row_reg, col_reg}<16'b1001000101111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000101111111) && ({row_reg, col_reg}<16'b1001000110000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001000110000011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001000110000100) && ({row_reg, col_reg}<16'b1001000110000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001000110000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000110001000) && ({row_reg, col_reg}<16'b1001000110001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001000110001010) && ({row_reg, col_reg}<16'b1001000110001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000110001101) && ({row_reg, col_reg}<16'b1001000110010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001000110010001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001000110010010) && ({row_reg, col_reg}<16'b1001000110010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001000110010100) && ({row_reg, col_reg}<16'b1001000110010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001000110010110) && ({row_reg, col_reg}<16'b1001000110100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001000110100011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001000110100100) && ({row_reg, col_reg}<16'b1001000110101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001000110101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000110101100) && ({row_reg, col_reg}<16'b1001000110110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001000110110001) && ({row_reg, col_reg}<16'b1001000110110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001000110110011) && ({row_reg, col_reg}<16'b1001000110110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001000110110101) && ({row_reg, col_reg}<16'b1001000110110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000110110111) && ({row_reg, col_reg}<16'b1001000110111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001000110111001) && ({row_reg, col_reg}<16'b1001000110111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001000111000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000111000001) && ({row_reg, col_reg}<16'b1001000111000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001000111000101)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==16'b1001000111000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001000111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000111001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001000111001001) && ({row_reg, col_reg}<16'b1001000111001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000111001100) && ({row_reg, col_reg}<16'b1001000111011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000111011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000111011010) && ({row_reg, col_reg}<16'b1001000111101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000111101000) && ({row_reg, col_reg}<16'b1001000111101010)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b1001000111101010) && ({row_reg, col_reg}<16'b1001001000001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001000001000) && ({row_reg, col_reg}<16'b1001001000001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001000001010) && ({row_reg, col_reg}<16'b1001001000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001000001101) && ({row_reg, col_reg}<16'b1001001000001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001001000001111) && ({row_reg, col_reg}<16'b1001001000010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001001000010011) && ({row_reg, col_reg}<16'b1001001000100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001000100101) && ({row_reg, col_reg}<16'b1001001000101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001000101001) && ({row_reg, col_reg}<16'b1001001000110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001000110010) && ({row_reg, col_reg}<16'b1001001000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001000110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001001000110110) && ({row_reg, col_reg}<16'b1001001000111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001000111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001001000111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001001000111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001000111011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1001001000111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001001000111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001001000111110) && ({row_reg, col_reg}<16'b1001001001000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001001001000000) && ({row_reg, col_reg}<16'b1001001001000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001001000010) && ({row_reg, col_reg}<16'b1001001001000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001001001000100) && ({row_reg, col_reg}<16'b1001001001000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001001000111) && ({row_reg, col_reg}<16'b1001001001001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001001001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001001001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001001001001011) && ({row_reg, col_reg}<16'b1001001001001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001001001101) && ({row_reg, col_reg}<16'b1001001001010000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001001001010000) && ({row_reg, col_reg}<16'b1001001001010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001001001010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001001010101) && ({row_reg, col_reg}<16'b1001001001011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001001001011010) && ({row_reg, col_reg}<16'b1001001001011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001001011100) && ({row_reg, col_reg}<16'b1001001001101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001001001101001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1001001001101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001001001101011) && ({row_reg, col_reg}<16'b1001001001101101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001001001101101) && ({row_reg, col_reg}<16'b1001001001111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001001001111101) && ({row_reg, col_reg}<16'b1001001010000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001010000010) && ({row_reg, col_reg}<16'b1001001010000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001001010000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001010000111) && ({row_reg, col_reg}<16'b1001001010001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001001010001001) && ({row_reg, col_reg}<16'b1001001010001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001010001011) && ({row_reg, col_reg}<16'b1001001010010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001001010010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001001010010001) && ({row_reg, col_reg}<16'b1001001010100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001001010100010) && ({row_reg, col_reg}<16'b1001001010100100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001001010100100) && ({row_reg, col_reg}<16'b1001001010101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001001010101001) && ({row_reg, col_reg}<16'b1001001010101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001010101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001001010101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001010101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001001010101110) && ({row_reg, col_reg}<16'b1001001010110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001010110001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001001010110010) && ({row_reg, col_reg}<16'b1001001010110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001001010110100) && ({row_reg, col_reg}<16'b1001001010110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001010110110) && ({row_reg, col_reg}<16'b1001001010111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001001010111000) && ({row_reg, col_reg}<16'b1001001010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001010111010) && ({row_reg, col_reg}<16'b1001001010111100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001001010111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001010111101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001001010111110) && ({row_reg, col_reg}<16'b1001001011000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001001011000000) && ({row_reg, col_reg}<16'b1001001011000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001011000010) && ({row_reg, col_reg}<16'b1001001011000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001011000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001001011000101) && ({row_reg, col_reg}<16'b1001001011000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001001011000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001011001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001001011001001) && ({row_reg, col_reg}<16'b1001001011001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001011001011) && ({row_reg, col_reg}<16'b1001001011010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001011010010) && ({row_reg, col_reg}<16'b1001001011010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001011010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001011010110) && ({row_reg, col_reg}<16'b1001001011011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001011011000) && ({row_reg, col_reg}<16'b1001001011100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001011100010) && ({row_reg, col_reg}<16'b1001001011100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001011100110) && ({row_reg, col_reg}<16'b1001001011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001011111001) && ({row_reg, col_reg}<16'b1001001011111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001011111100) && ({row_reg, col_reg}<16'b1001001011111111)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b1001001011111111) && ({row_reg, col_reg}<16'b1001001100001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001100001010) && ({row_reg, col_reg}<16'b1001001100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001100001101) && ({row_reg, col_reg}<16'b1001001100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001001100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001001100010010) && ({row_reg, col_reg}<16'b1001001100010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001100010110) && ({row_reg, col_reg}<16'b1001001100011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001100011000) && ({row_reg, col_reg}<16'b1001001100100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001100100110) && ({row_reg, col_reg}<16'b1001001100101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001100101000) && ({row_reg, col_reg}<16'b1001001100101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001100101110) && ({row_reg, col_reg}<16'b1001001100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001100110000) && ({row_reg, col_reg}<16'b1001001100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001100110011) && ({row_reg, col_reg}<16'b1001001100111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001100111010) && ({row_reg, col_reg}<16'b1001001100111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001001100111100) && ({row_reg, col_reg}<16'b1001001100111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001001100111111) && ({row_reg, col_reg}<16'b1001001101000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001101000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001001101000100) && ({row_reg, col_reg}<16'b1001001101000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001101000111) && ({row_reg, col_reg}<16'b1001001101001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001001101001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001001101001100)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b1001001101001101) && ({row_reg, col_reg}<16'b1001001101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001101001111) && ({row_reg, col_reg}<16'b1001001101010010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001001101010010) && ({row_reg, col_reg}<16'b1001001101010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001001101010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001101010110) && ({row_reg, col_reg}<16'b1001001101011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001001101011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001101011101) && ({row_reg, col_reg}<16'b1001001101100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001001101100011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001001101100100) && ({row_reg, col_reg}<16'b1001001101101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001001101101100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001001101101101) && ({row_reg, col_reg}<16'b1001001101111110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001001101111110) && ({row_reg, col_reg}<16'b1001001110000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001110000010) && ({row_reg, col_reg}<16'b1001001110000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001001110000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001110000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001001110000110) && ({row_reg, col_reg}<16'b1001001110001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001110001100) && ({row_reg, col_reg}<16'b1001001110001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001001110001111) && ({row_reg, col_reg}<16'b1001001110010001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001001110010001) && ({row_reg, col_reg}<16'b1001001110100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001001110100010) && ({row_reg, col_reg}<16'b1001001110100101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001001110100101) && ({row_reg, col_reg}<16'b1001001110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001001110100111) && ({row_reg, col_reg}<16'b1001001110101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001110101001) && ({row_reg, col_reg}<16'b1001001110101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001001110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001110101100) && ({row_reg, col_reg}<16'b1001001110101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001001110101110) && ({row_reg, col_reg}<16'b1001001110110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001110110000) && ({row_reg, col_reg}<16'b1001001110110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001001110110010)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==16'b1001001110110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001001110110100) && ({row_reg, col_reg}<16'b1001001110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001110111101) && ({row_reg, col_reg}<16'b1001001110111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001001110111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001111000000) && ({row_reg, col_reg}<16'b1001001111000010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001001111000010) && ({row_reg, col_reg}<16'b1001001111000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001111000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001001111000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001111000110) && ({row_reg, col_reg}<16'b1001001111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001111001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001001111001001) && ({row_reg, col_reg}<16'b1001001111001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001111001100) && ({row_reg, col_reg}<16'b1001001111010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001001111010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001111010100) && ({row_reg, col_reg}<16'b1001001111010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001001111010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001111011000) && ({row_reg, col_reg}<16'b1001001111100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001111100000) && ({row_reg, col_reg}<16'b1001001111100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001111100011) && ({row_reg, col_reg}<16'b1001001111101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001111101011) && ({row_reg, col_reg}<16'b1001001111101101)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b1001001111101101) && ({row_reg, col_reg}<16'b1001010000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010000000000) && ({row_reg, col_reg}<16'b1001010000000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001010000000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001010000001000) && ({row_reg, col_reg}<16'b1001010000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010000001101) && ({row_reg, col_reg}<16'b1001010000010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001010000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010000010001) && ({row_reg, col_reg}<16'b1001010000010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010000010110) && ({row_reg, col_reg}<16'b1001010000011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010000011000) && ({row_reg, col_reg}<16'b1001010000100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010000100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010000100101) && ({row_reg, col_reg}<16'b1001010000101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010000101001) && ({row_reg, col_reg}<16'b1001010000101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010000101100) && ({row_reg, col_reg}<16'b1001010000101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010000101110) && ({row_reg, col_reg}<16'b1001010000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010000110001) && ({row_reg, col_reg}<16'b1001010000110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010000110011) && ({row_reg, col_reg}<16'b1001010000111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001010000111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010000111101) && ({row_reg, col_reg}<16'b1001010000111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010000111111) && ({row_reg, col_reg}<16'b1001010001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001010001000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010001000111) && ({row_reg, col_reg}<16'b1001010001001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001010001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010001001100) && ({row_reg, col_reg}<16'b1001010001001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001010001001111) && ({row_reg, col_reg}<16'b1001010001010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010001010011) && ({row_reg, col_reg}<16'b1001010001010111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010001010111) && ({row_reg, col_reg}<16'b1001010001011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010001011011) && ({row_reg, col_reg}<16'b1001010001011101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001010001011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010001011110) && ({row_reg, col_reg}<16'b1001010001100100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001010001100100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001010001100101) && ({row_reg, col_reg}<16'b1001010001101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001010001101000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1001010001101001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001010001101010) && ({row_reg, col_reg}<16'b1001010001101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001010001101100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1001010001101101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001010001101110) && ({row_reg, col_reg}<16'b1001010001110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001010001110111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001010001111000) && ({row_reg, col_reg}<16'b1001010001111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001010001111111) && ({row_reg, col_reg}<16'b1001010010000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010010000010) && ({row_reg, col_reg}<16'b1001010010000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001010010000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010010000101) && ({row_reg, col_reg}<16'b1001010010000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001010010000111) && ({row_reg, col_reg}<16'b1001010010001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010010001001) && ({row_reg, col_reg}<16'b1001010010001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001010010001110) && ({row_reg, col_reg}<16'b1001010010010001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001010010010001) && ({row_reg, col_reg}<16'b1001010010011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001010010011000) && ({row_reg, col_reg}<16'b1001010010011010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001010010011010) && ({row_reg, col_reg}<16'b1001010010100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001010010100010) && ({row_reg, col_reg}<16'b1001010010100100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001010010100100) && ({row_reg, col_reg}<16'b1001010010100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001010010100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010010100111) && ({row_reg, col_reg}<16'b1001010010101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010010101001) && ({row_reg, col_reg}<16'b1001010010101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001010010101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001010010101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010010101110) && ({row_reg, col_reg}<16'b1001010010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001010010110101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1001010010110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001010010110111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001010010111000) && ({row_reg, col_reg}<16'b1001010010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010010111010) && ({row_reg, col_reg}<16'b1001010010111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001010010111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001010010111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010010111110) && ({row_reg, col_reg}<16'b1001010011000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010011000001) && ({row_reg, col_reg}<16'b1001010011000100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1001010011000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001010011000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001010011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001010011000111) && ({row_reg, col_reg}<16'b1001010011001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010011001100) && ({row_reg, col_reg}<16'b1001010011100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010011100000) && ({row_reg, col_reg}<16'b1001010011100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010011100011) && ({row_reg, col_reg}<16'b1001010011101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010011101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001010011101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010011101010) && ({row_reg, col_reg}<16'b1001010011101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010011101101) && ({row_reg, col_reg}<16'b1001010011111110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b1001010011111110) && ({row_reg, col_reg}<16'b1001010100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010100000101) && ({row_reg, col_reg}<16'b1001010100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010100000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001010100001000) && ({row_reg, col_reg}<16'b1001010100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010100001101) && ({row_reg, col_reg}<16'b1001010100001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001010100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001010100010000) && ({row_reg, col_reg}<16'b1001010100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010100010010) && ({row_reg, col_reg}<16'b1001010100100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010100100011) && ({row_reg, col_reg}<16'b1001010100100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010100100110) && ({row_reg, col_reg}<16'b1001010100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010100101001) && ({row_reg, col_reg}<16'b1001010100101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001010100101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010100101110) && ({row_reg, col_reg}<16'b1001010100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010100110100) && ({row_reg, col_reg}<16'b1001010100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010100110110) && ({row_reg, col_reg}<16'b1001010100111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001010100111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001010100111011) && ({row_reg, col_reg}<16'b1001010100111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001010100111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010100111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010100111111) && ({row_reg, col_reg}<16'b1001010101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001010101000100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001010101000101) && ({row_reg, col_reg}<16'b1001010101001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010101001000) && ({row_reg, col_reg}<16'b1001010101001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001010101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010101001100) && ({row_reg, col_reg}<16'b1001010101001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001010101001110) && ({row_reg, col_reg}<16'b1001010101010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001010101010011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001010101010100) && ({row_reg, col_reg}<16'b1001010101011000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010101011000) && ({row_reg, col_reg}<16'b1001010101011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010101011011) && ({row_reg, col_reg}<16'b1001010101011111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001010101011111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010101100000) && ({row_reg, col_reg}<16'b1001010101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010101100010) && ({row_reg, col_reg}<16'b1001010101101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001010101101000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001010101101001) && ({row_reg, col_reg}<16'b1001010101101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001010101101111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001010101110000) && ({row_reg, col_reg}<16'b1001010101110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001010101110110) && ({row_reg, col_reg}<16'b1001010101111000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001010101111000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001010101111001) && ({row_reg, col_reg}<16'b1001010101111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001010101111011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001010101111100) && ({row_reg, col_reg}<16'b1001010110000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001010110000010) && ({row_reg, col_reg}<16'b1001010110000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010110000100) && ({row_reg, col_reg}<16'b1001010110001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001010110001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001010110001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001010110001010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001010110001011) && ({row_reg, col_reg}<16'b1001010110001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001010110001111) && ({row_reg, col_reg}<16'b1001010110010001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001010110010001) && ({row_reg, col_reg}<16'b1001010110010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001010110010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001010110010111) && ({row_reg, col_reg}<16'b1001010110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001010110011010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001010110011011) && ({row_reg, col_reg}<16'b1001010110100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001010110100010) && ({row_reg, col_reg}<16'b1001010110100100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001010110100100) && ({row_reg, col_reg}<16'b1001010110100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001010110100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010110100111) && ({row_reg, col_reg}<16'b1001010110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010110101011) && ({row_reg, col_reg}<16'b1001010110101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001010110101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010110101110) && ({row_reg, col_reg}<16'b1001010110110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001010110110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001010110110111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001010110111000) && ({row_reg, col_reg}<16'b1001010110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010110111010) && ({row_reg, col_reg}<16'b1001010110111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001010110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001010110111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010110111111) && ({row_reg, col_reg}<16'b1001010111000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001010111000001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1001010111000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001010111000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010111000100) && ({row_reg, col_reg}<16'b1001010111000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001010111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001010111000111) && ({row_reg, col_reg}<16'b1001010111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010111001001) && ({row_reg, col_reg}<16'b1001010111100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010111100010) && ({row_reg, col_reg}<16'b1001010111100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001010111100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010111100111) && ({row_reg, col_reg}<16'b1001010111101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010111101101) && ({row_reg, col_reg}<16'b1001010111111101)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b1001010111111101) && ({row_reg, col_reg}<16'b1001011000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011000000110) && ({row_reg, col_reg}<16'b1001011000001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011000001000) && ({row_reg, col_reg}<16'b1001011000001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001011000001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001011000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011000001101) && ({row_reg, col_reg}<16'b1001011000001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001011000001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001011000010000) && ({row_reg, col_reg}<16'b1001011000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001011000010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011000010011) && ({row_reg, col_reg}<16'b1001011000011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001011000011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011000011011) && ({row_reg, col_reg}<16'b1001011000011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011000011110) && ({row_reg, col_reg}<16'b1001011000100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011000100001) && ({row_reg, col_reg}<16'b1001011000101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011000101001) && ({row_reg, col_reg}<16'b1001011000101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011000101100) && ({row_reg, col_reg}<16'b1001011000110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011000110011) && ({row_reg, col_reg}<16'b1001011000110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011000110111) && ({row_reg, col_reg}<16'b1001011000111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011000111001) && ({row_reg, col_reg}<16'b1001011000111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001011000111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001011000111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011000111111) && ({row_reg, col_reg}<16'b1001011001000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001011001000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001011001000010) && ({row_reg, col_reg}<16'b1001011001000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011001000100) && ({row_reg, col_reg}<16'b1001011001001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001011001001011) && ({row_reg, col_reg}<16'b1001011001001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001011001001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001011001001110) && ({row_reg, col_reg}<16'b1001011001010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011001010011) && ({row_reg, col_reg}<16'b1001011001010110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001011001010110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001011001010111) && ({row_reg, col_reg}<16'b1001011001011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011001011100) && ({row_reg, col_reg}<16'b1001011001100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001011001100000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011001100001) && ({row_reg, col_reg}<16'b1001011001100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011001100011) && ({row_reg, col_reg}<16'b1001011001100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001011001100101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001011001100110) && ({row_reg, col_reg}<16'b1001011001101011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1001011001101011) && ({row_reg, col_reg}<16'b1001011001101101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001011001101101) && ({row_reg, col_reg}<16'b1001011001110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001011001110000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001011001110001) && ({row_reg, col_reg}<16'b1001011001110011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001011001110011) && ({row_reg, col_reg}<16'b1001011001111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001011001111001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001011001111010) && ({row_reg, col_reg}<16'b1001011001111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1001011001111110) && ({row_reg, col_reg}<16'b1001011010000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001011010000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011010000100) && ({row_reg, col_reg}<16'b1001011010001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001011010001001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001011010001010) && ({row_reg, col_reg}<16'b1001011010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001011010001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001011010001101) && ({row_reg, col_reg}<16'b1001011010001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001011010001111) && ({row_reg, col_reg}<16'b1001011010010001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001011010010001) && ({row_reg, col_reg}<16'b1001011010010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001011010010101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001011010010110) && ({row_reg, col_reg}<16'b1001011010011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001011010011101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1001011010011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001011010011111) && ({row_reg, col_reg}<16'b1001011010100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001011010100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001011010100010) && ({row_reg, col_reg}<16'b1001011010100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001011010100101) && ({row_reg, col_reg}<16'b1001011010100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011010100111) && ({row_reg, col_reg}<16'b1001011010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011010101010) && ({row_reg, col_reg}<16'b1001011010101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011010101100) && ({row_reg, col_reg}<16'b1001011010101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001011010101111) && ({row_reg, col_reg}<16'b1001011010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001011010110011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001011010110100) && ({row_reg, col_reg}<16'b1001011010111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001011010111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001011010111010) && ({row_reg, col_reg}<16'b1001011010111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011010111100) && ({row_reg, col_reg}<16'b1001011010111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001011010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001011010111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011011000000) && ({row_reg, col_reg}<16'b1001011011000010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001011011000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011011000011) && ({row_reg, col_reg}<16'b1001011011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011011001001) && ({row_reg, col_reg}<16'b1001011011001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011011001111) && ({row_reg, col_reg}<16'b1001011011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011011010001) && ({row_reg, col_reg}<16'b1001011011011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011011011000) && ({row_reg, col_reg}<16'b1001011011101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011011101000) && ({row_reg, col_reg}<16'b1001011011101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011011101010) && ({row_reg, col_reg}<16'b1001011011101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011011101101) && ({row_reg, col_reg}<16'b1001011011110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011011110101) && ({row_reg, col_reg}<16'b1001011011111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011011111010) && ({row_reg, col_reg}<16'b1001011011111100)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b1001011011111100) && ({row_reg, col_reg}<16'b1001011100000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011100000111) && ({row_reg, col_reg}<16'b1001011100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011100001001) && ({row_reg, col_reg}<16'b1001011100001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001011100001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001011100001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001011100001110) && ({row_reg, col_reg}<16'b1001011100010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001011100010000) && ({row_reg, col_reg}<16'b1001011100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001011100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011100010011) && ({row_reg, col_reg}<16'b1001011100011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001011100011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011100011011) && ({row_reg, col_reg}<16'b1001011100011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011100011110) && ({row_reg, col_reg}<16'b1001011100100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011100100000) && ({row_reg, col_reg}<16'b1001011100101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011100101010) && ({row_reg, col_reg}<16'b1001011100101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011100101100) && ({row_reg, col_reg}<16'b1001011100110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011100110010) && ({row_reg, col_reg}<16'b1001011100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001011100110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001011100110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011100111000) && ({row_reg, col_reg}<16'b1001011100111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011100111011) && ({row_reg, col_reg}<16'b1001011100111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001011100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001011100111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001011101000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001011101000001) && ({row_reg, col_reg}<16'b1001011101000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001011101000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001011101000100) && ({row_reg, col_reg}<16'b1001011101000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011101000110) && ({row_reg, col_reg}<16'b1001011101001101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001011101001101) && ({row_reg, col_reg}<16'b1001011101010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001011101010000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1001011101010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011101010010) && ({row_reg, col_reg}<16'b1001011101010110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011101010110) && ({row_reg, col_reg}<16'b1001011101011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011101011001) && ({row_reg, col_reg}<16'b1001011101011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011101011100) && ({row_reg, col_reg}<16'b1001011101100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001011101100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011101100010) && ({row_reg, col_reg}<16'b1001011101100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001011101100100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001011101100101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001011101100110) && ({row_reg, col_reg}<16'b1001011101101010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001011101101010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001011101101011) && ({row_reg, col_reg}<16'b1001011101101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001011101101101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001011101101110) && ({row_reg, col_reg}<16'b1001011101110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1001011101110001) && ({row_reg, col_reg}<16'b1001011101110011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001011101110011) && ({row_reg, col_reg}<16'b1001011101111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001011101111110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001011101111111) && ({row_reg, col_reg}<16'b1001011110000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001011110000110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001011110000111) && ({row_reg, col_reg}<16'b1001011110001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001011110001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1001011110001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1001011110001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001011110001111) && ({row_reg, col_reg}<16'b1001011110010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001011110010011) && ({row_reg, col_reg}<16'b1001011110010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001011110010101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001011110010110) && ({row_reg, col_reg}<16'b1001011110011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001011110011000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1001011110011001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1001011110011010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001011110011011) && ({row_reg, col_reg}<16'b1001011110011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1001011110011110) && ({row_reg, col_reg}<16'b1001011110100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001011110100000) && ({row_reg, col_reg}<16'b1001011110100100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001011110100100) && ({row_reg, col_reg}<16'b1001011110100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011110100111) && ({row_reg, col_reg}<16'b1001011110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011110101001) && ({row_reg, col_reg}<16'b1001011110101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011110101011) && ({row_reg, col_reg}<16'b1001011110101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011110101101) && ({row_reg, col_reg}<16'b1001011110101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001011110101111) && ({row_reg, col_reg}<16'b1001011110110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001011110110001) && ({row_reg, col_reg}<16'b1001011110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001011110110011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001011110110100) && ({row_reg, col_reg}<16'b1001011110111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001011110111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001011110111010) && ({row_reg, col_reg}<16'b1001011111000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001011111000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011111000010) && ({row_reg, col_reg}<16'b1001011111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011111000101) && ({row_reg, col_reg}<16'b1001011111000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011111000111) && ({row_reg, col_reg}<16'b1001011111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011111001001) && ({row_reg, col_reg}<16'b1001011111001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011111001111) && ({row_reg, col_reg}<16'b1001011111010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011111010010) && ({row_reg, col_reg}<16'b1001011111010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011111010111) && ({row_reg, col_reg}<16'b1001011111100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001011111100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011111100101) && ({row_reg, col_reg}<16'b1001011111101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011111101000) && ({row_reg, col_reg}<16'b1001011111101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011111101010) && ({row_reg, col_reg}<16'b1001011111101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011111101101) && ({row_reg, col_reg}<16'b1001011111110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011111110101) && ({row_reg, col_reg}<16'b1001011111111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011111111010) && ({row_reg, col_reg}<16'b1001011111111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011111111100) && ({row_reg, col_reg}<16'b1001011111111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001011111111110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b1001011111111111) && ({row_reg, col_reg}<16'b1001100000000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100000000111) && ({row_reg, col_reg}<16'b1001100000001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100000001001) && ({row_reg, col_reg}<16'b1001100000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100000001100) && ({row_reg, col_reg}<16'b1001100000010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001100000010000) && ({row_reg, col_reg}<16'b1001100000011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100000011001) && ({row_reg, col_reg}<16'b1001100000011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100000011011) && ({row_reg, col_reg}<16'b1001100000011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100000011101) && ({row_reg, col_reg}<16'b1001100000011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001100000011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100000100000) && ({row_reg, col_reg}<16'b1001100000100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100000100011) && ({row_reg, col_reg}<16'b1001100000110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100000110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100000110111) && ({row_reg, col_reg}<16'b1001100000111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100000111011) && ({row_reg, col_reg}<16'b1001100000111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001100000111110) && ({row_reg, col_reg}<16'b1001100001000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100001000001) && ({row_reg, col_reg}<16'b1001100001000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001100001000100) && ({row_reg, col_reg}<16'b1001100001000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001100001000111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001100001001000) && ({row_reg, col_reg}<16'b1001100001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100001001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100001001100) && ({row_reg, col_reg}<16'b1001100001010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100001010000) && ({row_reg, col_reg}<16'b1001100001010010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001100001010010) && ({row_reg, col_reg}<16'b1001100001010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100001010100) && ({row_reg, col_reg}<16'b1001100001011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100001011000) && ({row_reg, col_reg}<16'b1001100001011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001100001011010) && ({row_reg, col_reg}<16'b1001100001100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100001100010) && ({row_reg, col_reg}<16'b1001100001100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001100001100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100001100101) && ({row_reg, col_reg}<16'b1001100001101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001100001101001) && ({row_reg, col_reg}<16'b1001100001101011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001100001101011) && ({row_reg, col_reg}<16'b1001100001101110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1001100001101110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1001100001101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001100001110000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001100001110001) && ({row_reg, col_reg}<16'b1001100001110011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001100001110011) && ({row_reg, col_reg}<16'b1001100001110110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1001100001110110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1001100001110111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001100001111000) && ({row_reg, col_reg}<16'b1001100001111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1001100001111010) && ({row_reg, col_reg}<16'b1001100001111101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1001100001111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1001100001111110) && ({row_reg, col_reg}<16'b1001100010000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001100010000100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001100010000101) && ({row_reg, col_reg}<16'b1001100010001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001100010001011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001100010001100) && ({row_reg, col_reg}<16'b1001100010001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001100010001110) && ({row_reg, col_reg}<16'b1001100010010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001100010010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001100010010001) && ({row_reg, col_reg}<16'b1001100010010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001100010010101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001100010010110) && ({row_reg, col_reg}<16'b1001100010011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001100010011000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1001100010011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001100010011010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001100010011011) && ({row_reg, col_reg}<16'b1001100010011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001100010011110) && ({row_reg, col_reg}<16'b1001100010100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001100010100000) && ({row_reg, col_reg}<16'b1001100010100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001100010100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100010100011) && ({row_reg, col_reg}<16'b1001100010100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100010100101) && ({row_reg, col_reg}<16'b1001100010101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100010101001) && ({row_reg, col_reg}<16'b1001100010101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100010101011) && ({row_reg, col_reg}<16'b1001100010101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100010101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001100010101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001100010110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001100010110001) && ({row_reg, col_reg}<16'b1001100010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100010110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001100010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001100010110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100010110111) && ({row_reg, col_reg}<16'b1001100010111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100010111011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001100010111100) && ({row_reg, col_reg}<16'b1001100011000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100011000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001100011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001100011000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100011000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001100011000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100011000101) && ({row_reg, col_reg}<16'b1001100011000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001100011000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100011001000) && ({row_reg, col_reg}<16'b1001100011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100011001010) && ({row_reg, col_reg}<16'b1001100011001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100011001100) && ({row_reg, col_reg}<16'b1001100011001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001100011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100011001111) && ({row_reg, col_reg}<16'b1001100011010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001100011010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100011010011) && ({row_reg, col_reg}<16'b1001100011011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100011011001) && ({row_reg, col_reg}<16'b1001100011100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100011100001) && ({row_reg, col_reg}<16'b1001100011100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100011100011) && ({row_reg, col_reg}<16'b1001100011101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100011101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100011101001) && ({row_reg, col_reg}<16'b1001100011101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100011101101) && ({row_reg, col_reg}<16'b1001100011110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100011110001) && ({row_reg, col_reg}<16'b1001100011110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100011110100) && ({row_reg, col_reg}<16'b1001100011111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100011111010) && ({row_reg, col_reg}<16'b1001100011111101)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b1001100011111101) && ({row_reg, col_reg}<16'b1001100100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100100000000) && ({row_reg, col_reg}<16'b1001100100001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100100001000) && ({row_reg, col_reg}<16'b1001100100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100100001100) && ({row_reg, col_reg}<16'b1001100100010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001100100010000) && ({row_reg, col_reg}<16'b1001100100010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100100010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100100010100) && ({row_reg, col_reg}<16'b1001100100011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100100011000) && ({row_reg, col_reg}<16'b1001100100011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100100011010) && ({row_reg, col_reg}<16'b1001100100011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100100011100) && ({row_reg, col_reg}<16'b1001100100011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100100011110) && ({row_reg, col_reg}<16'b1001100100100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100100100100) && ({row_reg, col_reg}<16'b1001100100101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100100101101) && ({row_reg, col_reg}<16'b1001100100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100100110001) && ({row_reg, col_reg}<16'b1001100100111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100100111001) && ({row_reg, col_reg}<16'b1001100100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100100111011) && ({row_reg, col_reg}<16'b1001100100111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100100111101) && ({row_reg, col_reg}<16'b1001100100111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001100100111111) && ({row_reg, col_reg}<16'b1001100101000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100101000100) && ({row_reg, col_reg}<16'b1001100101000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001100101000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001100101000111) && ({row_reg, col_reg}<16'b1001100101010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100101010010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001100101010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100101010100) && ({row_reg, col_reg}<16'b1001100101010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100101010111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001100101011000) && ({row_reg, col_reg}<16'b1001100101011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100101011011) && ({row_reg, col_reg}<16'b1001100101100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100101100110) && ({row_reg, col_reg}<16'b1001100101101000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1001100101101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100101101001) && ({row_reg, col_reg}<16'b1001100101101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001100101101100) && ({row_reg, col_reg}<16'b1001100101101110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001100101101110) && ({row_reg, col_reg}<16'b1001100101110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001100101110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001100101110011) && ({row_reg, col_reg}<16'b1001100101110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001100101110111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001100101111000) && ({row_reg, col_reg}<16'b1001100101111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1001100101111010) && ({row_reg, col_reg}<16'b1001100101111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001100101111101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001100101111110) && ({row_reg, col_reg}<16'b1001100110000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001100110000011) && ({row_reg, col_reg}<16'b1001100110001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1001100110001011) && ({row_reg, col_reg}<16'b1001100110001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001100110001101) && ({row_reg, col_reg}<16'b1001100110010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001100110010100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1001100110010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001100110010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001100110010111) && ({row_reg, col_reg}<16'b1001100110011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1001100110011001) && ({row_reg, col_reg}<16'b1001100110011011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001100110011011) && ({row_reg, col_reg}<16'b1001100110100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001100110100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100110100001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001100110100010) && ({row_reg, col_reg}<16'b1001100110101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100110101011) && ({row_reg, col_reg}<16'b1001100110101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100110101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001100110101110) && ({row_reg, col_reg}<16'b1001100110110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100110110001) && ({row_reg, col_reg}<16'b1001100110110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001100110110110) && ({row_reg, col_reg}<16'b1001100110111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100110111000) && ({row_reg, col_reg}<16'b1001100110111010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001100110111010) && ({row_reg, col_reg}<16'b1001100110111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001100111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001100111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100111000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001100111000011) && ({row_reg, col_reg}<16'b1001100111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100111000101) && ({row_reg, col_reg}<16'b1001100111001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100111001010) && ({row_reg, col_reg}<16'b1001100111001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100111001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100111001101) && ({row_reg, col_reg}<16'b1001100111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100111010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100111010010) && ({row_reg, col_reg}<16'b1001100111010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100111010100) && ({row_reg, col_reg}<16'b1001100111010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100111010110) && ({row_reg, col_reg}<16'b1001100111011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100111011001) && ({row_reg, col_reg}<16'b1001100111011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100111011101) && ({row_reg, col_reg}<16'b1001100111101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100111101001) && ({row_reg, col_reg}<16'b1001100111110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100111110001) && ({row_reg, col_reg}<16'b1001100111110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100111110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100111110111) && ({row_reg, col_reg}<16'b1001100111111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100111111101)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b1001100111111110) && ({row_reg, col_reg}<16'b1001101000001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101000001000) && ({row_reg, col_reg}<16'b1001101000001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101000001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101000001100) && ({row_reg, col_reg}<16'b1001101000010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001101000010000) && ({row_reg, col_reg}<16'b1001101000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101000010010) && ({row_reg, col_reg}<16'b1001101000010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101000010100) && ({row_reg, col_reg}<16'b1001101000011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101000011000) && ({row_reg, col_reg}<16'b1001101000011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101000011010) && ({row_reg, col_reg}<16'b1001101000100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101000100000) && ({row_reg, col_reg}<16'b1001101000101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101000101100) && ({row_reg, col_reg}<16'b1001101000101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001101000101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001101000101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001101000110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101000110001) && ({row_reg, col_reg}<16'b1001101000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001101000110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101000110101) && ({row_reg, col_reg}<16'b1001101000111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001101000111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101000111011) && ({row_reg, col_reg}<16'b1001101000111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101000111101) && ({row_reg, col_reg}<16'b1001101001000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001101001000000) && ({row_reg, col_reg}<16'b1001101001000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101001000100) && ({row_reg, col_reg}<16'b1001101001000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101001000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001101001000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101001001000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001101001001001) && ({row_reg, col_reg}<16'b1001101001010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101001010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101001010011) && ({row_reg, col_reg}<16'b1001101001010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101001010101) && ({row_reg, col_reg}<16'b1001101001010111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001101001010111) && ({row_reg, col_reg}<16'b1001101001011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101001011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001101001011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101001011100) && ({row_reg, col_reg}<16'b1001101001100000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001101001100000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1001101001100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101001100010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001101001100011) && ({row_reg, col_reg}<16'b1001101001101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001101001101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001101001101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101001101010) && ({row_reg, col_reg}<16'b1001101001101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001101001101100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1001101001101101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001101001101110) && ({row_reg, col_reg}<16'b1001101001110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001101001110010) && ({row_reg, col_reg}<16'b1001101001110100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1001101001110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001101001110101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1001101001110110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001101001110111) && ({row_reg, col_reg}<16'b1001101001111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001101001111010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001101001111011) && ({row_reg, col_reg}<16'b1001101001111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001101001111101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001101001111110) && ({row_reg, col_reg}<16'b1001101010000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001101010000011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001101010000100) && ({row_reg, col_reg}<16'b1001101010001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001101010001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001101010001101) && ({row_reg, col_reg}<16'b1001101010010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001101010010001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1001101010010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001101010010011) && ({row_reg, col_reg}<16'b1001101010010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1001101010010101) && ({row_reg, col_reg}<16'b1001101010010111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001101010010111) && ({row_reg, col_reg}<16'b1001101010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001101010011010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001101010011011) && ({row_reg, col_reg}<16'b1001101010011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001101010011101) && ({row_reg, col_reg}<16'b1001101010011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001101010011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101010100000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001101010100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001101010100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001101010100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001101010100100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1001101010100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101010100110) && ({row_reg, col_reg}<16'b1001101010101001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001101010101001) && ({row_reg, col_reg}<16'b1001101010101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001101010101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001101010101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001101010101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101010101111) && ({row_reg, col_reg}<16'b1001101010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101010110110) && ({row_reg, col_reg}<16'b1001101010111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001101010111001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1001101010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101010111011) && ({row_reg, col_reg}<16'b1001101010111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001101010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101010111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001101010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101011000000) && ({row_reg, col_reg}<16'b1001101011000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101011000100) && ({row_reg, col_reg}<16'b1001101011001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101011001101) && ({row_reg, col_reg}<16'b1001101011011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101011011010) && ({row_reg, col_reg}<16'b1001101011011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101011011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001101011011110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101011011111) && ({row_reg, col_reg}<16'b1001101011100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101011100001) && ({row_reg, col_reg}<16'b1001101011100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101011100101) && ({row_reg, col_reg}<16'b1001101011101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101011101000) && ({row_reg, col_reg}<16'b1001101011110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101011110100) && ({row_reg, col_reg}<16'b1001101011111111)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}==16'b1001101011111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001101100000000) && ({row_reg, col_reg}<16'b1001101100001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001101100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101100001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101100001100) && ({row_reg, col_reg}<16'b1001101100010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001101100010000) && ({row_reg, col_reg}<16'b1001101100011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101100011111) && ({row_reg, col_reg}<16'b1001101100101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101100101101) && ({row_reg, col_reg}<16'b1001101100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101100110000) && ({row_reg, col_reg}<16'b1001101100110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101100110010) && ({row_reg, col_reg}<16'b1001101100110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001101100110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001101100110111) && ({row_reg, col_reg}<16'b1001101101000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101101000001) && ({row_reg, col_reg}<16'b1001101101000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001101101000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101101000100) && ({row_reg, col_reg}<16'b1001101101000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101101000111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001101101001000) && ({row_reg, col_reg}<16'b1001101101001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101101001010) && ({row_reg, col_reg}<16'b1001101101001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001101101001100) && ({row_reg, col_reg}<16'b1001101101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101101001111) && ({row_reg, col_reg}<16'b1001101101010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001101101010010) && ({row_reg, col_reg}<16'b1001101101010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101101010100) && ({row_reg, col_reg}<16'b1001101101011000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001101101011000) && ({row_reg, col_reg}<16'b1001101101011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101101011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001101101011011) && ({row_reg, col_reg}<16'b1001101101011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101101011101) && ({row_reg, col_reg}<16'b1001101101100000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001101101100000) && ({row_reg, col_reg}<16'b1001101101100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101101100100) && ({row_reg, col_reg}<16'b1001101101100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101101100110) && ({row_reg, col_reg}<16'b1001101101101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101101101001) && ({row_reg, col_reg}<16'b1001101101101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001101101101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101101101100) && ({row_reg, col_reg}<16'b1001101101110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001101101110010) && ({row_reg, col_reg}<16'b1001101101110110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001101101110110) && ({row_reg, col_reg}<16'b1001101101111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1001101101111010) && ({row_reg, col_reg}<16'b1001101101111100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1001101101111100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1001101101111101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001101101111110) && ({row_reg, col_reg}<16'b1001101110000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001101110000011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1001101110000100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001101110000101) && ({row_reg, col_reg}<16'b1001101110000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1001101110000111) && ({row_reg, col_reg}<16'b1001101110001001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1001101110001001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1001101110001010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1001101110001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001101110001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001101110001101) && ({row_reg, col_reg}<16'b1001101110010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001101110010001) && ({row_reg, col_reg}<16'b1001101110010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001101110010011) && ({row_reg, col_reg}<16'b1001101110010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1001101110010101) && ({row_reg, col_reg}<16'b1001101110010111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001101110010111) && ({row_reg, col_reg}<16'b1001101110011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001101110011010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001101110011011) && ({row_reg, col_reg}<16'b1001101110011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001101110011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101110011111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101110100000) && ({row_reg, col_reg}<16'b1001101110100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001101110100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101110100011) && ({row_reg, col_reg}<16'b1001101110101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101110101010) && ({row_reg, col_reg}<16'b1001101110101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001101110101100) && ({row_reg, col_reg}<16'b1001101110101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101110101110) && ({row_reg, col_reg}<16'b1001101110110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101110110100) && ({row_reg, col_reg}<16'b1001101110110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001101110110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101110110111) && ({row_reg, col_reg}<16'b1001101110111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001101110111001) && ({row_reg, col_reg}<16'b1001101110111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101110111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001101110111100) && ({row_reg, col_reg}<16'b1001101110111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101110111111) && ({row_reg, col_reg}<16'b1001101111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001101111000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001101111000010) && ({row_reg, col_reg}<16'b1001101111000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101111000100) && ({row_reg, col_reg}<16'b1001101111001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101111001101) && ({row_reg, col_reg}<16'b1001101111010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001101111010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101111010001) && ({row_reg, col_reg}<16'b1001101111010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101111010111) && ({row_reg, col_reg}<16'b1001101111011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001101111011001) && ({row_reg, col_reg}<16'b1001101111101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101111101010) && ({row_reg, col_reg}<16'b1001101111110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101111110101) && ({row_reg, col_reg}<16'b1001101111111111)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}==16'b1001101111111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001110000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110000000001) && ({row_reg, col_reg}<16'b1001110000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110000001100) && ({row_reg, col_reg}<16'b1001110000010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001110000010000) && ({row_reg, col_reg}<16'b1001110000011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110000011110) && ({row_reg, col_reg}<16'b1001110000101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110000101110) && ({row_reg, col_reg}<16'b1001110000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110000110000) && ({row_reg, col_reg}<16'b1001110000110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110000110011) && ({row_reg, col_reg}<16'b1001110001000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110001000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001110001000011) && ({row_reg, col_reg}<16'b1001110001000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110001000111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001110001001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110001001001) && ({row_reg, col_reg}<16'b1001110001001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001110001001011) && ({row_reg, col_reg}<16'b1001110001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110001001111) && ({row_reg, col_reg}<16'b1001110001010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001110001010010) && ({row_reg, col_reg}<16'b1001110001010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110001010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001110001010101) && ({row_reg, col_reg}<16'b1001110001011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110001011000) && ({row_reg, col_reg}<16'b1001110001011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001110001011011) && ({row_reg, col_reg}<16'b1001110001011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110001011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001110001011110) && ({row_reg, col_reg}<16'b1001110001100001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001110001100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001110001100011) && ({row_reg, col_reg}<16'b1001110001100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110001100101) && ({row_reg, col_reg}<16'b1001110001101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001110001101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110001101001) && ({row_reg, col_reg}<16'b1001110001101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001110001101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001110001101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001110001101101) && ({row_reg, col_reg}<16'b1001110001110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110001110000) && ({row_reg, col_reg}<16'b1001110001110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001110001110011) && ({row_reg, col_reg}<16'b1001110001110110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001110001110110) && ({row_reg, col_reg}<16'b1001110001111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001110001111001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1001110001111010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001110001111011) && ({row_reg, col_reg}<16'b1001110001111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001110001111101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1001110001111110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001110001111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001110010000000) && ({row_reg, col_reg}<16'b1001110010000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001110010000011) && ({row_reg, col_reg}<16'b1001110010000111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001110010000111) && ({row_reg, col_reg}<16'b1001110010001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001110010001011) && ({row_reg, col_reg}<16'b1001110010010101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1001110010010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001110010010110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001110010010111) && ({row_reg, col_reg}<16'b1001110010011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1001110010011010) && ({row_reg, col_reg}<16'b1001110010011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001110010011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110010011101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001110010011110) && ({row_reg, col_reg}<16'b1001110010100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001110010100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001110010100100) && ({row_reg, col_reg}<16'b1001110010101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110010101001) && ({row_reg, col_reg}<16'b1001110010101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001110010101011) && ({row_reg, col_reg}<16'b1001110010101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110010101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001110010101110) && ({row_reg, col_reg}<16'b1001110010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110010110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001110010110011) && ({row_reg, col_reg}<16'b1001110010110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110010110110) && ({row_reg, col_reg}<16'b1001110010111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001110010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110010111001) && ({row_reg, col_reg}<16'b1001110010111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001110010111101) && ({row_reg, col_reg}<16'b1001110010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110010111111) && ({row_reg, col_reg}<16'b1001110011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110011000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001110011000010) && ({row_reg, col_reg}<16'b1001110011000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110011000100) && ({row_reg, col_reg}<16'b1001110011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110011001010) && ({row_reg, col_reg}<16'b1001110011001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110011001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110011001101) && ({row_reg, col_reg}<16'b1001110011010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110011010000) && ({row_reg, col_reg}<16'b1001110011010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110011010010) && ({row_reg, col_reg}<16'b1001110011010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110011010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110011010110) && ({row_reg, col_reg}<16'b1001110011101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110011101011) && ({row_reg, col_reg}<16'b1001110011110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110011110100) && ({row_reg, col_reg}<16'b1001110011110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110011110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110011111000) && ({row_reg, col_reg}<16'b1001110011111011)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b1001110011111011) && ({row_reg, col_reg}<16'b1001110100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110100000000) && ({row_reg, col_reg}<16'b1001110100001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110100001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001110100001001) && ({row_reg, col_reg}<16'b1001110100001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110100001100) && ({row_reg, col_reg}<16'b1001110100010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001110100010000) && ({row_reg, col_reg}<16'b1001110100011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110100011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001110100011001) && ({row_reg, col_reg}<16'b1001110100011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110100011101) && ({row_reg, col_reg}<16'b1001110100100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110100100011) && ({row_reg, col_reg}<16'b1001110100100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110100100110) && ({row_reg, col_reg}<16'b1001110100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110100101001) && ({row_reg, col_reg}<16'b1001110100101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110100101101) && ({row_reg, col_reg}<16'b1001110100101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110100101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110100110000) && ({row_reg, col_reg}<16'b1001110100110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110100110100) && ({row_reg, col_reg}<16'b1001110101000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110101000100) && ({row_reg, col_reg}<16'b1001110101000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001110101000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110101000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110101001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001110101001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110101001010) && ({row_reg, col_reg}<16'b1001110101010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001110101010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110101010001) && ({row_reg, col_reg}<16'b1001110101010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001110101010100) && ({row_reg, col_reg}<16'b1001110101010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110101010110) && ({row_reg, col_reg}<16'b1001110101011000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001110101011000) && ({row_reg, col_reg}<16'b1001110101011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110101011101) && ({row_reg, col_reg}<16'b1001110101011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001110101011111) && ({row_reg, col_reg}<16'b1001110101100001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001110101100001) && ({row_reg, col_reg}<16'b1001110101100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110101100110) && ({row_reg, col_reg}<16'b1001110101101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110101101000) && ({row_reg, col_reg}<16'b1001110101101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110101101011) && ({row_reg, col_reg}<16'b1001110101110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001110101110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110101110001) && ({row_reg, col_reg}<16'b1001110101110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001110101110110) && ({row_reg, col_reg}<16'b1001110101111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001110101111001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1001110101111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001110101111011) && ({row_reg, col_reg}<16'b1001110110000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001110110000000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001110110000001) && ({row_reg, col_reg}<16'b1001110110000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001110110000011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001110110000100) && ({row_reg, col_reg}<16'b1001110110000110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1001110110000110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001110110000111) && ({row_reg, col_reg}<16'b1001110110001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001110110001001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1001110110001010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001110110001011) && ({row_reg, col_reg}<16'b1001110110010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1001110110010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001110110010001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001110110010010) && ({row_reg, col_reg}<16'b1001110110010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001110110010110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001110110010111) && ({row_reg, col_reg}<16'b1001110110011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001110110011001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1001110110011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001110110011011) && ({row_reg, col_reg}<16'b1001110110011101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001110110011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110110011110) && ({row_reg, col_reg}<16'b1001110110100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110110100010) && ({row_reg, col_reg}<16'b1001110110100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110110100100) && ({row_reg, col_reg}<16'b1001110110100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001110110100111) && ({row_reg, col_reg}<16'b1001110110101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110110101001) && ({row_reg, col_reg}<16'b1001110110101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001110110101011) && ({row_reg, col_reg}<16'b1001110110101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110110101101) && ({row_reg, col_reg}<16'b1001110110110001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001110110110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001110110110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001110110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110110110100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001110110110101) && ({row_reg, col_reg}<16'b1001110110110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110110110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001110110111000)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b1001110110111001) && ({row_reg, col_reg}<16'b1001110110111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001110110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110110111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001110111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110111000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001110111000010) && ({row_reg, col_reg}<16'b1001110111000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110111000100) && ({row_reg, col_reg}<16'b1001110111001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110111001010) && ({row_reg, col_reg}<16'b1001110111001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110111001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110111001101) && ({row_reg, col_reg}<16'b1001110111001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110111001111) && ({row_reg, col_reg}<16'b1001110111010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110111010010) && ({row_reg, col_reg}<16'b1001110111010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110111010101) && ({row_reg, col_reg}<16'b1001110111010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110111010111) && ({row_reg, col_reg}<16'b1001110111101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110111101100) && ({row_reg, col_reg}<16'b1001110111110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110111110101) && ({row_reg, col_reg}<16'b1001110111110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110111110111) && ({row_reg, col_reg}<16'b1001110111111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110111111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110111111010) && ({row_reg, col_reg}<16'b1001110111111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110111111100) && ({row_reg, col_reg}<16'b1001110111111110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b1001110111111110) && ({row_reg, col_reg}<16'b1001111000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111000000000) && ({row_reg, col_reg}<16'b1001111000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111000001100) && ({row_reg, col_reg}<16'b1001111000010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001111000010000) && ({row_reg, col_reg}<16'b1001111000010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111000010100) && ({row_reg, col_reg}<16'b1001111000010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111000010110) && ({row_reg, col_reg}<16'b1001111000011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111000011011) && ({row_reg, col_reg}<16'b1001111000100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111000100011) && ({row_reg, col_reg}<16'b1001111000100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111000100110) && ({row_reg, col_reg}<16'b1001111000101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111000101001) && ({row_reg, col_reg}<16'b1001111000101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111000101101) && ({row_reg, col_reg}<16'b1001111001000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111001000000) && ({row_reg, col_reg}<16'b1001111001001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111001001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001111001001010) && ({row_reg, col_reg}<16'b1001111001010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111001010001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001111001010010) && ({row_reg, col_reg}<16'b1001111001011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111001011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001111001011011) && ({row_reg, col_reg}<16'b1001111001011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111001011111) && ({row_reg, col_reg}<16'b1001111001100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001111001100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111001100100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001111001100101) && ({row_reg, col_reg}<16'b1001111001100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111001100111) && ({row_reg, col_reg}<16'b1001111001101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111001101110) && ({row_reg, col_reg}<16'b1001111001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111001110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001111001110001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001111001110010) && ({row_reg, col_reg}<16'b1001111001110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001111001110110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1001111001110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001111001111000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1001111001111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001111001111010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001111001111011) && ({row_reg, col_reg}<16'b1001111010000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001111010000000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001111010000001) && ({row_reg, col_reg}<16'b1001111010000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001111010000100) && ({row_reg, col_reg}<16'b1001111010000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1001111010000110) && ({row_reg, col_reg}<16'b1001111010001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001111010001000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001111010001001) && ({row_reg, col_reg}<16'b1001111010001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001111010001011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001111010001100) && ({row_reg, col_reg}<16'b1001111010001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001111010001111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1001111010010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001111010010001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001111010010010) && ({row_reg, col_reg}<16'b1001111010010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001111010010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001111010010111) && ({row_reg, col_reg}<16'b1001111010011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001111010011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111010011011) && ({row_reg, col_reg}<16'b1001111010011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111010011110) && ({row_reg, col_reg}<16'b1001111010100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001111010100001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001111010100010) && ({row_reg, col_reg}<16'b1001111010101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111010101101) && ({row_reg, col_reg}<16'b1001111010101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001111010101111) && ({row_reg, col_reg}<16'b1001111010110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111010110111) && ({row_reg, col_reg}<16'b1001111010111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001111010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111010111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001111010111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111010111101) && ({row_reg, col_reg}<16'b1001111010111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111010111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001111011000000) && ({row_reg, col_reg}<16'b1001111011000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111011000100) && ({row_reg, col_reg}<16'b1001111011010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111011010010) && ({row_reg, col_reg}<16'b1001111011010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111011010101) && ({row_reg, col_reg}<16'b1001111011011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111011011001) && ({row_reg, col_reg}<16'b1001111011011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111011011100) && ({row_reg, col_reg}<16'b1001111011101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111011101001) && ({row_reg, col_reg}<16'b1001111011101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111011101101) && ({row_reg, col_reg}<16'b1001111011110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111011110101) && ({row_reg, col_reg}<16'b1001111011111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111011111000) && ({row_reg, col_reg}<16'b1001111011111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111011111100) && ({row_reg, col_reg}<16'b1001111011111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111011111110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b1001111011111111) && ({row_reg, col_reg}<16'b1001111100001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111100001011) && ({row_reg, col_reg}<16'b1001111100010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001111100010000) && ({row_reg, col_reg}<16'b1001111100010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111100010100) && ({row_reg, col_reg}<16'b1001111100010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111100010111) && ({row_reg, col_reg}<16'b1001111100011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111100011010) && ({row_reg, col_reg}<16'b1001111100100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001111100100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111100100101) && ({row_reg, col_reg}<16'b1001111100100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111100100111) && ({row_reg, col_reg}<16'b1001111100101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111100101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001111100101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111100101100) && ({row_reg, col_reg}<16'b1001111101000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111101000000) && ({row_reg, col_reg}<16'b1001111101001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111101001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001111101001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001111101001100) && ({row_reg, col_reg}<16'b1001111101010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111101010010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001111101010011) && ({row_reg, col_reg}<16'b1001111101011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111101011111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001111101100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111101100001)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==16'b1001111101100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001111101100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111101100100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1001111101100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001111101100110) && ({row_reg, col_reg}<16'b1001111101101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111101101000) && ({row_reg, col_reg}<16'b1001111101101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001111101101011) && ({row_reg, col_reg}<16'b1001111101101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111101101110) && ({row_reg, col_reg}<16'b1001111101110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111101110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001111101110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001111101110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111101110100) && ({row_reg, col_reg}<16'b1001111101110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001111101110110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1001111101110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001111101111000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1001111101111001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001111101111010) && ({row_reg, col_reg}<16'b1001111101111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001111101111111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001111110000000) && ({row_reg, col_reg}<16'b1001111110000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001111110000100) && ({row_reg, col_reg}<16'b1001111110000110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001111110000110) && ({row_reg, col_reg}<16'b1001111110001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001111110001001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1001111110001010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001111110001011) && ({row_reg, col_reg}<16'b1001111110001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001111110001111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1001111110010000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1001111110010001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001111110010010) && ({row_reg, col_reg}<16'b1001111110010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001111110010100) && ({row_reg, col_reg}<16'b1001111110010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001111110010110) && ({row_reg, col_reg}<16'b1001111110011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001111110011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111110011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111110011011) && ({row_reg, col_reg}<16'b1001111110011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111110011101) && ({row_reg, col_reg}<16'b1001111110011111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111110011111) && ({row_reg, col_reg}<16'b1001111110100001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1001111110100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001111110100010) && ({row_reg, col_reg}<16'b1001111110110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111110110111) && ({row_reg, col_reg}<16'b1001111110111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001111110111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111110111100) && ({row_reg, col_reg}<16'b1001111110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111110111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001111110111111) && ({row_reg, col_reg}<16'b1001111111000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111111000011) && ({row_reg, col_reg}<16'b1001111111010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111111010100) && ({row_reg, col_reg}<16'b1001111111010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111111010111) && ({row_reg, col_reg}<16'b1001111111011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001111111011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111111011011) && ({row_reg, col_reg}<16'b1001111111011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111111011101) && ({row_reg, col_reg}<16'b1001111111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111111011111) && ({row_reg, col_reg}<16'b1001111111101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111111101001) && ({row_reg, col_reg}<16'b1001111111101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111111101100) && ({row_reg, col_reg}<16'b1001111111110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001111111110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111111110111) && ({row_reg, col_reg}<16'b1001111111111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001111111111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111111111101) && ({row_reg, col_reg}<16'b1001111111111111)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b1001111111111111) && ({row_reg, col_reg}<=16'b1001111111111111)) color_data = 12'b000100010000;
	end
endmodule