module enemy_rom
	(
		input wire clk,
		input wire [6:0] row,
		input wire [5:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [6:0] row_reg;
	reg [5:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin
		if(({row_reg, col_reg}>=13'b0000000000000) && ({row_reg, col_reg}<13'b0000000010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0000000010001)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0000000010010)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0000000010011)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0000000010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0000000010101) && ({row_reg, col_reg}<13'b0000000010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000000010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=13'b0000000011000) && ({row_reg, col_reg}<13'b0000000011101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0000000011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=13'b0000000011110) && ({row_reg, col_reg}<13'b0000000100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000000100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0000000100010) && ({row_reg, col_reg}<13'b0000000100101)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0000000100101)) color_data = 12'b010010010011;

		if(({row_reg, col_reg}>=13'b0000000100110) && ({row_reg, col_reg}<13'b0000001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0000001010000)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0000001010001)) color_data = 12'b001101110010;
		if(({row_reg, col_reg}>=13'b0000001010010) && ({row_reg, col_reg}<13'b0000001010101)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0000001010101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0000001010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000001010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0000001011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000001011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=13'b0000001011010) && ({row_reg, col_reg}<13'b0000001011100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=13'b0000001011100) && ({row_reg, col_reg}<13'b0000001011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0000001011111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000001100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0000001100001)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0000001100010)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0000001100011)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}>=13'b0000001100100) && ({row_reg, col_reg}<13'b0000001100110)) color_data = 12'b001101110010;
		if(({row_reg, col_reg}==13'b0000001100110)) color_data = 12'b001110000010;

		if(({row_reg, col_reg}>=13'b0000001100111) && ({row_reg, col_reg}<13'b0000010010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0000010010000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000010010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0000010010010)) color_data = 12'b001001010001;
		if(({row_reg, col_reg}==13'b0000010010011)) color_data = 12'b001101110010;
		if(({row_reg, col_reg}==13'b0000010010100)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0000010010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0000010010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000010010111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=13'b0000010011000) && ({row_reg, col_reg}<13'b0000010011100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=13'b0000010011100) && ({row_reg, col_reg}<13'b0000010011111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0000010011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0000010100000) && ({row_reg, col_reg}<13'b0000010100010)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0000010100010)) color_data = 12'b001101110010;
		if(({row_reg, col_reg}==13'b0000010100011)) color_data = 12'b001001010001;
		if(({row_reg, col_reg}>=13'b0000010100100) && ({row_reg, col_reg}<13'b0000010100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000010100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0000010100111)) color_data = 12'b001101110010;

		if(({row_reg, col_reg}>=13'b0000010101000) && ({row_reg, col_reg}<13'b0000011001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0000011001000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0000011001001) && ({row_reg, col_reg}<13'b0000011001011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b0000011001011) && ({row_reg, col_reg}<13'b0000011001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0000011001101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0000011001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0000011001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0000011010000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0000011010001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=13'b0000011010010) && ({row_reg, col_reg}<13'b0000011010100)) color_data = 12'b001001010001;
		if(({row_reg, col_reg}==13'b0000011010100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=13'b0000011010101) && ({row_reg, col_reg}<13'b0000011010111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=13'b0000011010111) && ({row_reg, col_reg}<13'b0000011011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=13'b0000011011001) && ({row_reg, col_reg}<13'b0000011011011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0000011011011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0000011011100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0000011011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0000011011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0000011011111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000011100000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0000011100001)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b0000011100010)) color_data = 12'b001001010001;
		if(({row_reg, col_reg}==13'b0000011100011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=13'b0000011100100) && ({row_reg, col_reg}<13'b0000011100110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0000011100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0000011100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0000011101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=13'b0000011101010) && ({row_reg, col_reg}<13'b0000011101100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0000011101100)) color_data = 12'b011001100110;

		if(({row_reg, col_reg}>=13'b0000011101101) && ({row_reg, col_reg}<13'b0000100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0000100000110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0000100000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0000100001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0000100001001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0000100001010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0000100001011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=13'b0000100001100) && ({row_reg, col_reg}<13'b0000100001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0000100001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0000100001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0000100010000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=13'b0000100010001) && ({row_reg, col_reg}<13'b0000100010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000100010011)) color_data = 12'b001001010001;
		if(({row_reg, col_reg}==13'b0000100010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0000100010101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0000100010110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0000100010111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=13'b0000100011000) && ({row_reg, col_reg}<13'b0000100011011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=13'b0000100011011) && ({row_reg, col_reg}<13'b0000100011101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0000100011101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0000100011111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0000100100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000100100001)) color_data = 12'b001001010001;
		if(({row_reg, col_reg}>=13'b0000100100010) && ({row_reg, col_reg}<13'b0000100100100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=13'b0000100100100) && ({row_reg, col_reg}<13'b0000100100110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0000100100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0000100100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000100101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=13'b0000100101001) && ({row_reg, col_reg}<13'b0000100101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0000100101011) && ({row_reg, col_reg}<13'b0000100101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0000100101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0000100101110)) color_data = 12'b010101010101;

		if(({row_reg, col_reg}>=13'b0000100101111) && ({row_reg, col_reg}<13'b0000101000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0000101000101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0000101000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0000101000111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0000101001000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0000101001001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0000101001010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0000101001011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0000101001101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0000101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0000101001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0000101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0000101010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000101010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0000101010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0000101010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0000101010101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0000101010110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0000101010111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0000101011000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0000101011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0000101011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=13'b0000101011011) && ({row_reg, col_reg}<13'b0000101011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0000101011101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0000101011110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0000101011111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0000101100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0000101100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0000101100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0000101100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0000101100100) && ({row_reg, col_reg}<13'b0000101100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=13'b0000101100110) && ({row_reg, col_reg}<13'b0000101101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0000101101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0000101101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0000101101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=13'b0000101101011) && ({row_reg, col_reg}<13'b0000101101101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0000101101101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0000101101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0000101101111)) color_data = 12'b010101010101;

		if(({row_reg, col_reg}>=13'b0000101110000) && ({row_reg, col_reg}<13'b0000110000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0000110000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0000110000101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0000110000110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000110000111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=13'b0000110001000) && ({row_reg, col_reg}<13'b0000110001010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0000110001010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0000110001011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0000110001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0000110001101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b0000110001110) && ({row_reg, col_reg}<13'b0000110010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0000110010000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0000110010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000110010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0000110010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000110010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0000110010101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000110010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=13'b0000110010111) && ({row_reg, col_reg}<13'b0000110011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0000110011001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=13'b0000110011010) && ({row_reg, col_reg}<13'b0000110100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000110100000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0000110100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0000110100010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0000110100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0000110100100) && ({row_reg, col_reg}<13'b0000110100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0000110100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000110100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0000110101000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0000110101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0000110101010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=13'b0000110101011) && ({row_reg, col_reg}<13'b0000110101101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0000110101101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0000110101110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0000110101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0000110110000)) color_data = 12'b010001000100;

		if(({row_reg, col_reg}>=13'b0000110110001) && ({row_reg, col_reg}<13'b0000111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0000111000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0000111000101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0000111000110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000111000111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0000111001000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0000111001001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0000111001010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0000111001011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000111001100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0000111001101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0000111001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0000111001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0000111010000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0000111010001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0000111010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0000111010011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0000111010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0000111010101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000111010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=13'b0000111010111) && ({row_reg, col_reg}<13'b0000111011001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=13'b0000111011001) && ({row_reg, col_reg}<13'b0000111011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=13'b0000111011011) && ({row_reg, col_reg}<13'b0000111011101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000111011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0000111011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0000111011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0000111100000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0000111100001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0000111100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0000111100011) && ({row_reg, col_reg}<13'b0000111100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0000111100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=13'b0000111100111) && ({row_reg, col_reg}<13'b0000111101001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0000111101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0000111101010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=13'b0000111101011) && ({row_reg, col_reg}<13'b0000111101101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0000111101101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0000111101110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0000111101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0000111110000)) color_data = 12'b001100110011;

		if(({row_reg, col_reg}>=13'b0000111110001) && ({row_reg, col_reg}<13'b0001000000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0001000000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001000000101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001000000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=13'b0001000000111) && ({row_reg, col_reg}<13'b0001000001001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001000001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0001000001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001000001011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001000001100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001000001101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0001000001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001000001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0001000010000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001000010001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001000010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0001000010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001000010100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0001000010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0001000010110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0001000010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001000011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0001000011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0001000011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0001000011011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0001000011100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0001000011101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=13'b0001000011110) && ({row_reg, col_reg}<13'b0001000100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0001000100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001000100001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0001000100010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001000100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0001000100100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001000100101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0001000100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=13'b0001000100111) && ({row_reg, col_reg}<13'b0001000101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001000101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001000101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=13'b0001000101011) && ({row_reg, col_reg}<13'b0001000101101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0001000101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0001000101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001000101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001000110000)) color_data = 12'b001100110011;

		if(({row_reg, col_reg}>=13'b0001000110001) && ({row_reg, col_reg}<13'b0001001000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0001001000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001001000101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001001000110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001001000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0001001001000) && ({row_reg, col_reg}<13'b0001001001011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001001001011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001001001100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0001001001101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001001001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0001001001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001001010000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001001010001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0001001010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0001001010011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001001010100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0001001010101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0001001010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001001010111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001001011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001001011001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001001011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0001001011011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0001001011100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0001001011101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0001001011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0001001011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001001100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0001001100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001001100010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001001100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0001001100100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0001001100101) && ({row_reg, col_reg}<13'b0001001100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0001001100111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0001001101000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0001001101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0001001101010) && ({row_reg, col_reg}<13'b0001001101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0001001101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001001101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001001110000)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=13'b0001001110001) && ({row_reg, col_reg}<13'b0001010000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0001010000011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0001010000100) && ({row_reg, col_reg}<13'b0001010000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0001010000110) && ({row_reg, col_reg}<13'b0001010001100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001010001100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0001010001101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001010001110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0001010001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001010010000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001010010001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0001010010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001010010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0001010010100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001010010101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=13'b0001010010110) && ({row_reg, col_reg}<13'b0001010011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0001010011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0001010011001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001010011010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0001010011011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0001010011100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b0001010011101) && ({row_reg, col_reg}<13'b0001010011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0001010011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0001010100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0001010100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001010100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001010100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001010100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001010100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001010100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0001010100111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0001010101000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0001010101001) && ({row_reg, col_reg}<13'b0001010101100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001010101100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b0001010101101) && ({row_reg, col_reg}<13'b0001010101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001010101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0001010110000)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}==13'b0001010110001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0001011000000) && ({row_reg, col_reg}<13'b0001011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0001011000011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001011000100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001011000101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0001011000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0001011000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0001011001000) && ({row_reg, col_reg}<13'b0001011001011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0001011001011) && ({row_reg, col_reg}<13'b0001011001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001011001101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001011001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0001011001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0001011010000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001011010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001011010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0001011010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0001011010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001011010101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0001011010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0001011010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0001011011000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001011011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0001011011010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0001011011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0001011011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0001011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0001011011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001011011111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001011100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0001011100001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0001011100010) && ({row_reg, col_reg}<13'b0001011100100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001011100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0001011100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0001011100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0001011100111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0001011101000) && ({row_reg, col_reg}<13'b0001011101110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001011101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0001011101111) && ({row_reg, col_reg}<13'b0001011110001)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}==13'b0001011110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0001100000000) && ({row_reg, col_reg}<13'b0001100000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0001100000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0001100000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0001100000101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0001100000110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001100000111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001100001000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001100001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001100001010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0001100001011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001100001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0001100001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0001100001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0001100001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001100010000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0001100010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0001100010011) && ({row_reg, col_reg}<13'b0001100010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0001100010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0001100010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001100010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0001100011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001100011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0001100011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001100011011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001100011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0001100011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0001100011110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001100011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0001100100000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001100100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001100100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001100100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001100100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001100100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001100100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=13'b0001100100111) && ({row_reg, col_reg}<13'b0001100101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001100101001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0001100101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001100101011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0001100101100) && ({row_reg, col_reg}<13'b0001100101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001100101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001100110000)) color_data = 12'b011001100110;

		if(({row_reg, col_reg}==13'b0001100110001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0001101000000) && ({row_reg, col_reg}<13'b0001101000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0001101000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001101000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001101000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0001101000110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=13'b0001101000111) && ({row_reg, col_reg}<13'b0001101001001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0001101001001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0001101001010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0001101001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=13'b0001101001100) && ({row_reg, col_reg}<13'b0001101001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0001101001110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0001101001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0001101010000) && ({row_reg, col_reg}<13'b0001101010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001101010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0001101010011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001101010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001101010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0001101010110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0001101010111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0001101011000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=13'b0001101011001) && ({row_reg, col_reg}<13'b0001101011011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001101011011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001101011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0001101011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001101011110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0001101011111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0001101100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001101100001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0001101100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001101100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0001101100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0001101100101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001101100110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0001101100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001101101000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0001101101001) && ({row_reg, col_reg}<13'b0001101101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0001101101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001101101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0001101110000)) color_data = 12'b011001100110;

		if(({row_reg, col_reg}==13'b0001101110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b0001110000000) && ({row_reg, col_reg}<13'b0001110000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0001110000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001110000101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001110000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0001110000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0001110001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001110001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0001110001010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0001110001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0001110001100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0001110001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0001110001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0001110001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0001110010000) && ({row_reg, col_reg}<13'b0001110010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001110010010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001110010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0001110010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0001110010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0001110010110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0001110010111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0001110011000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0001110011001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0001110011010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0001110011011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001110011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=13'b0001110011101) && ({row_reg, col_reg}<13'b0001110011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0001110011111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001110100000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0001110100001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0001110100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0001110100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001110100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0001110100101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0001110100110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=13'b0001110100111) && ({row_reg, col_reg}<13'b0001110101001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0001110101001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0001110101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0001110101011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=13'b0001110101100) && ({row_reg, col_reg}<13'b0001110101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0001110101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0001110101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001110110000)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=13'b0001110110001) && ({row_reg, col_reg}<13'b0001111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0001111000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0001111000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001111000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0001111000111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0001111001000) && ({row_reg, col_reg}<13'b0001111001010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0001111001010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0001111001011) && ({row_reg, col_reg}<13'b0001111001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0001111001101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0001111001110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001111001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b0001111010000) && ({row_reg, col_reg}<13'b0001111010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001111010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001111010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001111010101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0001111010110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0001111010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001111011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0001111011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0001111011010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=13'b0001111011011) && ({row_reg, col_reg}<13'b0001111011110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0001111011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b0001111011111) && ({row_reg, col_reg}<13'b0001111100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001111100010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0001111100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001111100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0001111100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001111100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0001111100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0001111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0001111101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0001111101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0001111101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0001111101100) && ({row_reg, col_reg}<13'b0001111101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0001111101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001111101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0001111110000)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=13'b0001111110001) && ({row_reg, col_reg}<13'b0010000000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0010000000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=13'b0010000000101) && ({row_reg, col_reg}<13'b0010000000111)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=13'b0010000000111) && ({row_reg, col_reg}<13'b0010000001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0010000001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0010000001010) && ({row_reg, col_reg}<13'b0010000001100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0010000001100) && ({row_reg, col_reg}<13'b0010000001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0010000001111) && ({row_reg, col_reg}<13'b0010000010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0010000010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0010000010100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0010000010101) && ({row_reg, col_reg}<13'b0010000010111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=13'b0010000010111) && ({row_reg, col_reg}<13'b0010000011001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0010000011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0010000011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0010000011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0010000011100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0010000011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0010000011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=13'b0010000011111) && ({row_reg, col_reg}<13'b0010000100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0010000100001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0010000100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0010000100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0010000100100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==13'b0010000100101)) color_data = 12'b000100110000;
		if(({row_reg, col_reg}>=13'b0010000100110) && ({row_reg, col_reg}<13'b0010000101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0010000101000) && ({row_reg, col_reg}<13'b0010000101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0010000101010) && ({row_reg, col_reg}<13'b0010000101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0010000101100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==13'b0010000101101)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==13'b0010000101110)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==13'b0010000101111)) color_data = 12'b001100110010;

		if(({row_reg, col_reg}>=13'b0010000110000) && ({row_reg, col_reg}<13'b0010001000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0010001000100)) color_data = 12'b001101110010;
		if(({row_reg, col_reg}>=13'b0010001000101) && ({row_reg, col_reg}<13'b0010001000111)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}>=13'b0010001000111) && ({row_reg, col_reg}<13'b0010001001001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==13'b0010001001001)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==13'b0010001001010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==13'b0010001001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=13'b0010001001100) && ({row_reg, col_reg}<13'b0010001001111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==13'b0010001001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0010001010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0010001010001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0010001010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0010001010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0010001010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0010001010101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0010001010110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0010001010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0010001011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0010001011001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0010001011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0010001011011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b0010001011100) && ({row_reg, col_reg}<13'b0010001011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0010001011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0010001011111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0010001100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0010001100001) && ({row_reg, col_reg}<13'b0010001100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0010001100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0010001100101)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=13'b0010001100110) && ({row_reg, col_reg}<13'b0010001101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==13'b0010001101000)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b0010001101001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==13'b0010001101010)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==13'b0010001101011)) color_data = 12'b001101110010;
		if(({row_reg, col_reg}==13'b0010001101100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==13'b0010001101101)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b0010001101110)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0010001101111)) color_data = 12'b001101110010;

		if(({row_reg, col_reg}>=13'b0010001110000) && ({row_reg, col_reg}<13'b0010010000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0010010000011)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==13'b0010010000100)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0010010000101)) color_data = 12'b011011010101;
		if(({row_reg, col_reg}==13'b0010010000110)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0010010000111)) color_data = 12'b010111000101;
		if(({row_reg, col_reg}>=13'b0010010001000) && ({row_reg, col_reg}<13'b0010010001010)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b0010010001010)) color_data = 12'b001101110010;
		if(({row_reg, col_reg}==13'b0010010001011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==13'b0010010001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=13'b0010010001101) && ({row_reg, col_reg}<13'b0010010001111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==13'b0010010001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0010010010000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0010010010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0010010010010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0010010010011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0010010010100) && ({row_reg, col_reg}<13'b0010010010110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0010010010110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=13'b0010010010111) && ({row_reg, col_reg}<13'b0010010011001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0010010011001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0010010011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0010010011011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0010010011100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0010010011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0010010011110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0010010011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0010010100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0010010100001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0010010100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0010010100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0010010100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0010010100101)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}>=13'b0010010100110) && ({row_reg, col_reg}<13'b0010010101000)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0010010101000)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0010010101001)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0010010101010)) color_data = 12'b011011100110;
		if(({row_reg, col_reg}==13'b0010010101011)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0010010101100)) color_data = 12'b011011100110;
		if(({row_reg, col_reg}==13'b0010010101101)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}>=13'b0010010101110) && ({row_reg, col_reg}<13'b0010010110000)) color_data = 12'b001110000010;

		if(({row_reg, col_reg}>=13'b0010010110000) && ({row_reg, col_reg}<13'b0010011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0010011000011)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==13'b0010011000100)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0010011000101)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0010011000110)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0010011000111)) color_data = 12'b011011100110;
		if(({row_reg, col_reg}==13'b0010011001000)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b0010011001001)) color_data = 12'b010110110100;
		if(({row_reg, col_reg}==13'b0010011001010)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==13'b0010011001011)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b0010011001100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==13'b0010011001101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==13'b0010011001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0010011001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0010011010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0010011010001) && ({row_reg, col_reg}<13'b0010011010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0010011010011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0010011010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0010011010101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0010011010110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0010011010111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=13'b0010011011000) && ({row_reg, col_reg}<13'b0010011011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0010011011010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0010011011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0010011011100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0010011011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0010011011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0010011011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0010011100000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0010011100001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0010011100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0010011100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0010011100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0010011100101)) color_data = 12'b001101110010;
		if(({row_reg, col_reg}==13'b0010011100110)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0010011100111)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0010011101000)) color_data = 12'b010110110100;
		if(({row_reg, col_reg}==13'b0010011101001)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0010011101010)) color_data = 12'b011111110110;
		if(({row_reg, col_reg}==13'b0010011101011)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0010011101100)) color_data = 12'b011011100110;
		if(({row_reg, col_reg}==13'b0010011101101)) color_data = 12'b001101110010;
		if(({row_reg, col_reg}==13'b0010011101110)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0010011101111)) color_data = 12'b001001100010;

		if(({row_reg, col_reg}>=13'b0010011110000) && ({row_reg, col_reg}<13'b0010100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0010100000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0010100000010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0010100000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0010100000100)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0010100000101)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}>=13'b0010100000110) && ({row_reg, col_reg}<13'b0010100001000)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0010100001000)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0010100001001)) color_data = 12'b010110110100;
		if(({row_reg, col_reg}==13'b0010100001010)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==13'b0010100001011)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0010100001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0010100001101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==13'b0010100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0010100001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0010100010000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0010100010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0010100010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0010100010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0010100010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0010100010101) && ({row_reg, col_reg}<13'b0010100010111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0010100010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0010100011000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0010100011001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0010100011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0010100011011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0010100011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0010100011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0010100011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0010100011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0010100100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0010100100001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0010100100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0010100100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0010100100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0010100100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==13'b0010100100110)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0010100100111)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0010100101000)) color_data = 12'b010110110100;
		if(({row_reg, col_reg}==13'b0010100101001)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0010100101010)) color_data = 12'b011011100110;
		if(({row_reg, col_reg}==13'b0010100101011)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0010100101100)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}>=13'b0010100101101) && ({row_reg, col_reg}<13'b0010100101111)) color_data = 12'b001101110010;
		if(({row_reg, col_reg}==13'b0010100101111)) color_data = 12'b001100110010;

		if(({row_reg, col_reg}>=13'b0010100110000) && ({row_reg, col_reg}<13'b0010101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0010101000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0010101000010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0010101000011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=13'b0010101000100) && ({row_reg, col_reg}<13'b0010101000110)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==13'b0010101000110)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0010101000111)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b0010101001000)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0010101001001)) color_data = 12'b001101110010;
		if(({row_reg, col_reg}==13'b0010101001010)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0010101001011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==13'b0010101001100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=13'b0010101001101) && ({row_reg, col_reg}<13'b0010101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0010101001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0010101010000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0010101010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0010101010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0010101010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0010101010101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0010101010110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0010101010111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0010101011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0010101011001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0010101011010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0010101011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0010101011100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0010101011101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0010101011110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0010101011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0010101100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0010101100001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0010101100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0010101100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0010101100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0010101100101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==13'b0010101100110)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0010101100111)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b0010101101000)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0010101101001)) color_data = 12'b001101110010;
		if(({row_reg, col_reg}==13'b0010101101010)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0010101101011)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0010101101100)) color_data = 12'b001101110010;
		if(({row_reg, col_reg}==13'b0010101101101)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b0010101101110)) color_data = 12'b001101110010;

		if(({row_reg, col_reg}>=13'b0010101101111) && ({row_reg, col_reg}<13'b0010110000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0010110000000) && ({row_reg, col_reg}<13'b0010110000010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==13'b0010110000010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0010110000011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==13'b0010110000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0010110000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==13'b0010110000110)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b0010110000111)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==13'b0010110001000)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0010110001001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==13'b0010110001010)) color_data = 12'b001101110010;
		if(({row_reg, col_reg}==13'b0010110001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0010110001100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=13'b0010110001101) && ({row_reg, col_reg}<13'b0010110010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0010110010000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0010110010001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b0010110010010) && ({row_reg, col_reg}<13'b0010110010100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0010110010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0010110010101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0010110010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0010110010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0010110011000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b0010110011001) && ({row_reg, col_reg}<13'b0010110011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0010110011011) && ({row_reg, col_reg}<13'b0010110011101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0010110011101) && ({row_reg, col_reg}<13'b0010110011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0010110011111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0010110100000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0010110100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0010110100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0010110100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0010110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==13'b0010110100101)) color_data = 12'b000100110000;
		if(({row_reg, col_reg}>=13'b0010110100110) && ({row_reg, col_reg}<13'b0010110101000)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b0010110101000)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0010110101001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==13'b0010110101010)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0010110101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==13'b0010110101100)) color_data = 12'b001101110010;
		if(({row_reg, col_reg}==13'b0010110101101)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b0010110101110)) color_data = 12'b001100110010;

		if(({row_reg, col_reg}>=13'b0010110101111) && ({row_reg, col_reg}<13'b0010111000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0010111000000)) color_data = 12'b110110110100;
		if(({row_reg, col_reg}==13'b0010111000001)) color_data = 12'b110010010010;
		if(({row_reg, col_reg}==13'b0010111000010)) color_data = 12'b011001110101;
		if(({row_reg, col_reg}==13'b0010111000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0010111000100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==13'b0010111000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0010111000110)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==13'b0010111000111)) color_data = 12'b001101110010;
		if(({row_reg, col_reg}==13'b0010111001000)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==13'b0010111001001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==13'b0010111001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0010111001011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=13'b0010111001100) && ({row_reg, col_reg}<13'b0010111010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0010111010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0010111010001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0010111010010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0010111010011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0010111010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0010111010101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0010111010110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0010111010111) && ({row_reg, col_reg}<13'b0010111011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0010111011001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0010111011010) && ({row_reg, col_reg}<13'b0010111011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0010111011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0010111011101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0010111011110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0010111011111) && ({row_reg, col_reg}<13'b0010111100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0010111100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0010111100010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0010111100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0010111100100) && ({row_reg, col_reg}<13'b0010111100110)) color_data = 12'b000100110000;
		if(({row_reg, col_reg}==13'b0010111100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==13'b0010111100111)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==13'b0010111101000)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b0010111101001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==13'b0010111101010)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}>=13'b0010111101011) && ({row_reg, col_reg}<13'b0010111101110)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==13'b0010111101110)) color_data = 12'b001001010001;

		if(({row_reg, col_reg}>=13'b0010111101111) && ({row_reg, col_reg}<13'b0011000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0011000000000)) color_data = 12'b111111110110;
		if(({row_reg, col_reg}==13'b0011000000001)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==13'b0011000000010)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0011000000011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0011000000100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=13'b0011000000101) && ({row_reg, col_reg}<13'b0011000000111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=13'b0011000000111) && ({row_reg, col_reg}<13'b0011000001001)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==13'b0011000001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=13'b0011000001010) && ({row_reg, col_reg}<13'b0011000001100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=13'b0011000001100) && ({row_reg, col_reg}<13'b0011000010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0011000010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0011000010010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0011000010011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0011000010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0011000010101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0011000010110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0011000010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0011000011000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b0011000011001) && ({row_reg, col_reg}<13'b0011000011011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0011000011011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0011000011100) && ({row_reg, col_reg}<13'b0011000011110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0011000011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0011000011111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0011000100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0011000100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0011000100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0011000100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0011000100100) && ({row_reg, col_reg}<13'b0011000100110)) color_data = 12'b000100110000;
		if(({row_reg, col_reg}==13'b0011000100110)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==13'b0011000100111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==13'b0011000101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==13'b0011000101001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==13'b0011000101010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==13'b0011000101011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=13'b0011000101100) && ({row_reg, col_reg}<13'b0011000101110)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=13'b0011000101110) && ({row_reg, col_reg}<13'b0011000110000)) color_data = 12'b001001010001;

		if(({row_reg, col_reg}>=13'b0011000110000) && ({row_reg, col_reg}<13'b0011001000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0011001000000) && ({row_reg, col_reg}<13'b0011001000010)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==13'b0011001000010)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0011001000011)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0011001000100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0011001000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0011001000110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0011001000111) && ({row_reg, col_reg}<13'b0011001001010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==13'b0011001001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b0011001001011) && ({row_reg, col_reg}<13'b0011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0011001010001) && ({row_reg, col_reg}<13'b0011001010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0011001010110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0011001010111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0011001011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0011001011001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0011001011010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0011001011011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0011001011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0011001011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0011001011110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0011001011111) && ({row_reg, col_reg}<13'b0011001100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0011001100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b0011001100010) && ({row_reg, col_reg}<13'b0011001100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0011001100100) && ({row_reg, col_reg}<13'b0011001100110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==13'b0011001100110)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==13'b0011001100111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==13'b0011001101000)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==13'b0011001101001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==13'b0011001101010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0011001101011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0011001101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0011001101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0011001101110)) color_data = 12'b001001010001;
		if(({row_reg, col_reg}>=13'b0011001101111) && ({row_reg, col_reg}<13'b0011001110001)) color_data = 12'b001101110010;

		if(({row_reg, col_reg}==13'b0011001110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0011010000000)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b0011010000001)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0011010000010)) color_data = 12'b110010010010;
		if(({row_reg, col_reg}==13'b0011010000011)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0011010000100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0011010000101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0011010000110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0011010000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0011010001000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==13'b0011010001001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0011010001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0011010001011) && ({row_reg, col_reg}<13'b0011010010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0011010010000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0011010010001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0011010010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0011010010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0011010010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0011010010101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0011010010110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0011010010111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0011010011000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0011010011001) && ({row_reg, col_reg}<13'b0011010011011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0011010011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0011010011100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0011010011101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0011010011110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0011010011111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0011010100000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0011010100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0011010100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0011010100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b0011010100100) && ({row_reg, col_reg}<13'b0011010100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0011010100110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0011010100111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0011010101000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0011010101001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0011010101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0011010101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0011010101100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0011010101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0011010101110)) color_data = 12'b001001010001;
		if(({row_reg, col_reg}==13'b0011010101111)) color_data = 12'b001101110010;
		if(({row_reg, col_reg}==13'b0011010110000)) color_data = 12'b001110000010;

		if(({row_reg, col_reg}==13'b0011010110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0011011000000)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b0011011000001)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0011011000010)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0011011000011)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0011011000100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0011011000101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0011011000110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0011011000111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0011011001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0011011001001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0011011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b0011011001011) && ({row_reg, col_reg}<13'b0011011001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0011011001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0011011010000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0011011010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0011011010010) && ({row_reg, col_reg}<13'b0011011010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0011011010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0011011010101) && ({row_reg, col_reg}<13'b0011011010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0011011010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0011011011000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0011011011001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0011011011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0011011011011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b0011011011100) && ({row_reg, col_reg}<13'b0011011011110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0011011011110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0011011011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b0011011100000) && ({row_reg, col_reg}<13'b0011011100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0011011100010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0011011100011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0011011100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0011011100101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0011011100110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0011011100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0011011101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0011011101001) && ({row_reg, col_reg}<13'b0011011101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0011011101011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0011011101100) && ({row_reg, col_reg}<13'b0011011101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0011011101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0011011101111)) color_data = 12'b001001010001;
		if(({row_reg, col_reg}==13'b0011011110000)) color_data = 12'b010010010011;

		if(({row_reg, col_reg}==13'b0011011110001)) color_data = 12'b001101110010;
		if(({row_reg, col_reg}==13'b0011100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0011100000001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b0011100000010) && ({row_reg, col_reg}<13'b0011100000100)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0011100000100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=13'b0011100000101) && ({row_reg, col_reg}<13'b0011100000111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0011100000111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0011100001000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0011100001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0011100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b0011100001011) && ({row_reg, col_reg}<13'b0011100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0011100001110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0011100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b0011100010000) && ({row_reg, col_reg}<13'b0011100010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0011100010011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0011100010100) && ({row_reg, col_reg}<13'b0011100010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0011100010110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0011100010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0011100011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0011100011001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=13'b0011100011010) && ({row_reg, col_reg}<13'b0011100011100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0011100011100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0011100011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0011100011110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0011100011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0011100100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0011100100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0011100100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0011100100011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0011100100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0011100100101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0011100100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0011100100111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0011100101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0011100101001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0011100101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0011100101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0011100101100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0011100101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0011100101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0011100101111)) color_data = 12'b001001010001;

		if(({row_reg, col_reg}>=13'b0011100110000) && ({row_reg, col_reg}<13'b0011101000000)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0011101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0011101000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0011101000010)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==13'b0011101000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==13'b0011101000100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0011101000101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0011101000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0011101000111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0011101001000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0011101001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0011101001010) && ({row_reg, col_reg}<13'b0011101001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0011101001110) && ({row_reg, col_reg}<13'b0011101010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0011101010101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0011101010110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0011101010111) && ({row_reg, col_reg}<13'b0011101011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0011101011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=13'b0011101011010) && ({row_reg, col_reg}<13'b0011101011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0011101011100) && ({row_reg, col_reg}<13'b0011101011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0011101011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0011101011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0011101100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0011101100001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0011101100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0011101100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0011101100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0011101100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0011101100110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0011101100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0011101101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0011101101001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0011101101010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0011101101011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0011101101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0011101101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0011101101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0011101101111)) color_data = 12'b001001010001;
		if(({row_reg, col_reg}==13'b0011101110000)) color_data = 12'b001101110010;

		if(({row_reg, col_reg}==13'b0011101110001)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0011110000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0011110000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0011110000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0011110000011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0011110000100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0011110000101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0011110000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0011110000111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0011110001000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0011110001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0011110001010) && ({row_reg, col_reg}<13'b0011110001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0011110001101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0011110001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0011110001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0011110010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0011110010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0011110010010) && ({row_reg, col_reg}<13'b0011110010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0011110010100) && ({row_reg, col_reg}<13'b0011110010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0011110010111) && ({row_reg, col_reg}<13'b0011110011001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b0011110011001) && ({row_reg, col_reg}<13'b0011110011011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0011110011011) && ({row_reg, col_reg}<13'b0011110011101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0011110011101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0011110011110) && ({row_reg, col_reg}<13'b0011110100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0011110100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0011110100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0011110100010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=13'b0011110100011) && ({row_reg, col_reg}<13'b0011110100101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0011110100101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0011110100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0011110100111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0011110101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0011110101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0011110101010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0011110101011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0011110101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0011110101101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0011110101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0011110101111)) color_data = 12'b001001010001;
		if(({row_reg, col_reg}==13'b0011110110000)) color_data = 12'b001110000010;

		if(({row_reg, col_reg}==13'b0011110110001)) color_data = 12'b001101110010;
		if(({row_reg, col_reg}==13'b0011111000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0011111000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0011111000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0011111000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0011111000100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0011111000101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0011111000110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0011111000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0011111001000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0011111001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0011111001010) && ({row_reg, col_reg}<13'b0011111001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0011111001100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0011111001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0011111001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0011111001111) && ({row_reg, col_reg}<13'b0011111010001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0011111010001) && ({row_reg, col_reg}<13'b0011111010011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0011111010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0011111010100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0011111010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0011111010110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0011111010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0011111011000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0011111011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0011111011010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0011111011011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0011111011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0011111011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0011111011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0011111011111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==13'b0011111100000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==13'b0011111100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==13'b0011111100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0011111100011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==13'b0011111100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==13'b0011111100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==13'b0011111100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==13'b0011111100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==13'b0011111101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==13'b0011111101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0011111101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0011111101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0011111101100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0011111101101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0011111101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0011111101111)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0011111110000)) color_data = 12'b010010010011;

		if(({row_reg, col_reg}==13'b0011111110001)) color_data = 12'b001101110010;
		if(({row_reg, col_reg}==13'b0100000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0100000000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0100000000010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0100000000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0100000000100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0100000000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==13'b0100000000110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0100000000111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b0100000001000) && ({row_reg, col_reg}<13'b0100000001010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0100000001010) && ({row_reg, col_reg}<13'b0100000001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0100000001100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0100000001101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0100000001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0100000001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0100000010000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0100000010001) && ({row_reg, col_reg}<13'b0100000010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0100000010011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0100000010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0100000010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0100000010110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0100000010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0100000011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=13'b0100000011001) && ({row_reg, col_reg}<13'b0100000011011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0100000011011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0100000011100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0100000011101)) color_data = 12'b101000110011;
		if(({row_reg, col_reg}==13'b0100000011110)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}>=13'b0100000011111) && ({row_reg, col_reg}<13'b0100000100001)) color_data = 12'b101000110011;
		if(({row_reg, col_reg}>=13'b0100000100001) && ({row_reg, col_reg}<13'b0100000100100)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==13'b0100000100100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==13'b0100000100101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==13'b0100000100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0100000100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==13'b0100000101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=13'b0100000101001) && ({row_reg, col_reg}<13'b0100000101011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0100000101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0100000101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0100000101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0100000101110)) color_data = 12'b001001010001;
		if(({row_reg, col_reg}>=13'b0100000101111) && ({row_reg, col_reg}<13'b0100000110001)) color_data = 12'b010010010011;

		if(({row_reg, col_reg}==13'b0100000110001)) color_data = 12'b001001010001;
		if(({row_reg, col_reg}==13'b0100001000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0100001000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0100001000010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0100001000011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0100001000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0100001000101)) color_data = 12'b110010010010;
		if(({row_reg, col_reg}>=13'b0100001000110) && ({row_reg, col_reg}<13'b0100001001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0100001001001) && ({row_reg, col_reg}<13'b0100001001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0100001001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0100001001100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0100001001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=13'b0100001001110) && ({row_reg, col_reg}<13'b0100001010000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0100001010000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0100001010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0100001010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0100001010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0100001010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0100001010101) && ({row_reg, col_reg}<13'b0100001010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0100001010111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0100001011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=13'b0100001011001) && ({row_reg, col_reg}<13'b0100001011011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0100001011011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0100001011100)) color_data = 12'b101101010101;
		if(({row_reg, col_reg}>=13'b0100001011101) && ({row_reg, col_reg}<13'b0100001011111)) color_data = 12'b101000110011;
		if(({row_reg, col_reg}>=13'b0100001011111) && ({row_reg, col_reg}<13'b0100001100001)) color_data = 12'b101101010101;
		if(({row_reg, col_reg}==13'b0100001100001)) color_data = 12'b101000110011;
		if(({row_reg, col_reg}==13'b0100001100010)) color_data = 12'b101101010101;
		if(({row_reg, col_reg}>=13'b0100001100011) && ({row_reg, col_reg}<13'b0100001100101)) color_data = 12'b101000110011;
		if(({row_reg, col_reg}==13'b0100001100101)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==13'b0100001100110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==13'b0100001100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==13'b0100001101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0100001101001) && ({row_reg, col_reg}<13'b0100001101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0100001101011) && ({row_reg, col_reg}<13'b0100001101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0100001101101)) color_data = 12'b001001010001;
		if(({row_reg, col_reg}>=13'b0100001101110) && ({row_reg, col_reg}<13'b0100001110000)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0100001110000)) color_data = 12'b001101110010;

		if(({row_reg, col_reg}==13'b0100001110001)) color_data = 12'b001001010001;
		if(({row_reg, col_reg}==13'b0100010000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0100010000001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0100010000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0100010000011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0100010000100)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==13'b0100010000101)) color_data = 12'b111111110100;
		if(({row_reg, col_reg}==13'b0100010000110)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}>=13'b0100010000111) && ({row_reg, col_reg}<13'b0100010001001)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}>=13'b0100010001001) && ({row_reg, col_reg}<13'b0100010001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0100010001011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0100010001100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0100010001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0100010001110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0100010001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0100010010000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0100010010001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0100010010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0100010010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0100010010100) && ({row_reg, col_reg}<13'b0100010010110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0100010010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0100010010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0100010011000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0100010011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0100010011010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0100010011011)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==13'b0100010011100)) color_data = 12'b110001100110;
		if(({row_reg, col_reg}==13'b0100010011101)) color_data = 12'b101000110011;
		if(({row_reg, col_reg}==13'b0100010011110)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==13'b0100010011111)) color_data = 12'b101000110011;
		if(({row_reg, col_reg}==13'b0100010100000)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==13'b0100010100001)) color_data = 12'b101000110011;
		if(({row_reg, col_reg}==13'b0100010100010)) color_data = 12'b101101000100;
		if(({row_reg, col_reg}>=13'b0100010100011) && ({row_reg, col_reg}<13'b0100010100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==13'b0100010100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0100010100110)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==13'b0100010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0100010101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0100010101001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0100010101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0100010101011) && ({row_reg, col_reg}<13'b0100010101101)) color_data = 12'b001001010001;
		if(({row_reg, col_reg}>=13'b0100010101101) && ({row_reg, col_reg}<13'b0100010110000)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0100010110000)) color_data = 12'b001001010001;

		if(({row_reg, col_reg}>=13'b0100010110001) && ({row_reg, col_reg}<13'b0100011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0100011000001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0100011000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0100011000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0100011000100)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==13'b0100011000101)) color_data = 12'b110110110100;
		if(({row_reg, col_reg}==13'b0100011000110)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0100011000111)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}>=13'b0100011001000) && ({row_reg, col_reg}<13'b0100011001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0100011001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0100011001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0100011001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=13'b0100011001101) && ({row_reg, col_reg}<13'b0100011001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0100011001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0100011010000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0100011010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0100011010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0100011010011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0100011010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0100011010101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0100011010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0100011010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0100011011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0100011011001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0100011011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0100011011011)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==13'b0100011011100)) color_data = 12'b101101000100;
		if(({row_reg, col_reg}>=13'b0100011011101) && ({row_reg, col_reg}<13'b0100011011111)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==13'b0100011011111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==13'b0100011100000)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==13'b0100011100001)) color_data = 12'b101101010101;
		if(({row_reg, col_reg}==13'b0100011100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==13'b0100011100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==13'b0100011100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==13'b0100011100101)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==13'b0100011100110)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==13'b0100011100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0100011101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0100011101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0100011101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0100011101011)) color_data = 12'b001101110010;
		if(({row_reg, col_reg}>=13'b0100011101100) && ({row_reg, col_reg}<13'b0100011101111)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0100011101111)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b0100011110000)) color_data = 12'b001001010001;

		if(({row_reg, col_reg}>=13'b0100011110001) && ({row_reg, col_reg}<13'b0100100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0100100000001) && ({row_reg, col_reg}<13'b0100100000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0100100000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0100100000100)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0100100000101)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}>=13'b0100100000110) && ({row_reg, col_reg}<13'b0100100001000)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b0100100001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0100100001001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0100100001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0100100001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0100100001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0100100001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0100100001110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0100100001111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0100100010000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0100100010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0100100010010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0100100010011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0100100010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0100100010101) && ({row_reg, col_reg}<13'b0100100011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b0100100011000) && ({row_reg, col_reg}<13'b0100100011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0100100011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==13'b0100100011100)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}>=13'b0100100011101) && ({row_reg, col_reg}<13'b0100100100000)) color_data = 12'b101000110011;
		if(({row_reg, col_reg}==13'b0100100100000)) color_data = 12'b101101010101;
		if(({row_reg, col_reg}==13'b0100100100001)) color_data = 12'b101000110011;
		if(({row_reg, col_reg}>=13'b0100100100010) && ({row_reg, col_reg}<13'b0100100100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==13'b0100100100100)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==13'b0100100100101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==13'b0100100100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0100100100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==13'b0100100101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0100100101001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0100100101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0100100101011)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}>=13'b0100100101100) && ({row_reg, col_reg}<13'b0100100101110)) color_data = 12'b001101110010;
		if(({row_reg, col_reg}==13'b0100100101110)) color_data = 12'b001001010001;
		if(({row_reg, col_reg}==13'b0100100101111)) color_data = 12'b000101000001;

		if(({row_reg, col_reg}>=13'b0100100110000) && ({row_reg, col_reg}<13'b0100101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0100101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0100101000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0100101000011)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0100101000100)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0100101000101)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0100101000110)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}>=13'b0100101000111) && ({row_reg, col_reg}<13'b0100101001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0100101001001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0100101001010) && ({row_reg, col_reg}<13'b0100101001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0100101001100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0100101001101)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0100101001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0100101001111) && ({row_reg, col_reg}<13'b0100101010001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0100101010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0100101010010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0100101010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0100101010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0100101010101)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b0100101010110)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0100101010111)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}>=13'b0100101011000) && ({row_reg, col_reg}<13'b0100101011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0100101011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0100101011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==13'b0100101011101)) color_data = 12'b110001100110;
		if(({row_reg, col_reg}==13'b0100101011110)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}==13'b0100101011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0100101100000)) color_data = 12'b110001100110;
		if(({row_reg, col_reg}==13'b0100101100001)) color_data = 12'b101101000100;
		if(({row_reg, col_reg}==13'b0100101100010)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==13'b0100101100011)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==13'b0100101100100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0100101100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==13'b0100101100110)) color_data = 12'b101000110011;
		if(({row_reg, col_reg}==13'b0100101100111)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==13'b0100101101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0100101101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0100101101010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b0100101101011) && ({row_reg, col_reg}<13'b0100101101101)) color_data = 12'b001001010001;
		if(({row_reg, col_reg}==13'b0100101101101)) color_data = 12'b000100110000;

		if(({row_reg, col_reg}>=13'b0100101101110) && ({row_reg, col_reg}<13'b0100110000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0100110000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0100110000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0100110000011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0100110000100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0100110000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0100110000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0100110000111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0100110001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0100110001001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0100110001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0100110001011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0100110001100)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0100110001101)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0100110001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0100110001111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0100110010000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0100110010001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0100110010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0100110010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0100110010100)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0100110010101)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0100110010110)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0100110010111)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}>=13'b0100110011000) && ({row_reg, col_reg}<13'b0100110011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0100110011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0100110011100)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==13'b0100110011101)) color_data = 12'b101101010101;
		if(({row_reg, col_reg}>=13'b0100110011110) && ({row_reg, col_reg}<13'b0100110100000)) color_data = 12'b110001100110;
		if(({row_reg, col_reg}==13'b0100110100000)) color_data = 12'b101101000100;
		if(({row_reg, col_reg}==13'b0100110100001)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==13'b0100110100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==13'b0100110100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=13'b0100110100100) && ({row_reg, col_reg}<13'b0100110100110)) color_data = 12'b000100110000;
		if(({row_reg, col_reg}==13'b0100110100110)) color_data = 12'b101101000100;
		if(({row_reg, col_reg}==13'b0100110100111)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==13'b0100110101000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0100110101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0100110101010)) color_data = 12'b010001000100;

		if(({row_reg, col_reg}>=13'b0100110101011) && ({row_reg, col_reg}<13'b0100111000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0100111000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0100111000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0100111000011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0100111000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0100111000101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0100111000110) && ({row_reg, col_reg}<13'b0100111001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0100111001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0100111001001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0100111001010) && ({row_reg, col_reg}<13'b0100111001100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0100111001100)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0100111001101)) color_data = 12'b110010010010;
		if(({row_reg, col_reg}==13'b0100111001110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0100111001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0100111010000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0100111010001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0100111010010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==13'b0100111010011)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0100111010100)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0100111010101)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0100111010110)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}>=13'b0100111010111) && ({row_reg, col_reg}<13'b0100111011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0100111011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==13'b0100111011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0100111011101)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==13'b0100111011110)) color_data = 12'b101000110011;
		if(({row_reg, col_reg}==13'b0100111011111)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==13'b0100111100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==13'b0100111100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==13'b0100111100010)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0100111100011)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0100111100100)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0100111100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0100111100110)) color_data = 12'b101000110011;
		if(({row_reg, col_reg}==13'b0100111100111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==13'b0100111101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0100111101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0100111101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0100111101011)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=13'b0100111101100) && ({row_reg, col_reg}<13'b0101000000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0101000000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0101000000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0101000000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0101000000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0101000000101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0101000000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0101000000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0101000001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0101000001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0101000001010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0101000001011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0101000001100)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0101000001101)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0101000001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0101000001111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0101000010000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0101000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0101000010010)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0101000010011)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0101000010100)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0101000010101)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}>=13'b0101000010110) && ({row_reg, col_reg}<13'b0101000011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0101000011011)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0101000011100)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}>=13'b0101000011101) && ({row_reg, col_reg}<13'b0101000100000)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==13'b0101000100000)) color_data = 12'b110010010010;
		if(({row_reg, col_reg}==13'b0101000100001)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0101000100010)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0101000100011)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0101000100100)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0101000100101)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==13'b0101000100110)) color_data = 12'b101000110011;
		if(({row_reg, col_reg}==13'b0101000100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=13'b0101000101000) && ({row_reg, col_reg}<13'b0101000101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0101000101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0101000101011)) color_data = 12'b100110011001;

		if(({row_reg, col_reg}>=13'b0101000101100) && ({row_reg, col_reg}<13'b0101001000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0101001000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b0101001000011) && ({row_reg, col_reg}<13'b0101001000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0101001000101) && ({row_reg, col_reg}<13'b0101001000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0101001000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0101001001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0101001001001) && ({row_reg, col_reg}<13'b0101001001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0101001001011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0101001001100)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0101001001101)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0101001001110)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}>=13'b0101001001111) && ({row_reg, col_reg}<13'b0101001010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0101001010010)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0101001010011)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0101001010100)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}>=13'b0101001010101) && ({row_reg, col_reg}<13'b0101001011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0101001011011)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0101001011100)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0101001011101)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0101001011110)) color_data = 12'b110010010010;
		if(({row_reg, col_reg}==13'b0101001011111)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}>=13'b0101001100000) && ({row_reg, col_reg}<13'b0101001100011)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0101001100011)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0101001100100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==13'b0101001100101)) color_data = 12'b101000110011;
		if(({row_reg, col_reg}==13'b0101001100110)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==13'b0101001100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==13'b0101001101000)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0101001101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0101001101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0101001101011)) color_data = 12'b011101110111;

		if(({row_reg, col_reg}>=13'b0101001101100) && ({row_reg, col_reg}<13'b0101010000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0101010000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0101010000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0101010000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b0101010000110) && ({row_reg, col_reg}<13'b0101010001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0101010001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0101010001001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0101010001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0101010001011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0101010001100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=13'b0101010001101) && ({row_reg, col_reg}<13'b0101010001111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0101010001111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0101010010000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0101010010001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0101010010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0101010010011)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}>=13'b0101010010100) && ({row_reg, col_reg}<13'b0101010011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0101010011011)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0101010011100)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0101010011101)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==13'b0101010011110)) color_data = 12'b111111110110;
		if(({row_reg, col_reg}==13'b0101010011111)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=13'b0101010100000) && ({row_reg, col_reg}<13'b0101010100010)) color_data = 12'b110110110100;
		if(({row_reg, col_reg}==13'b0101010100010)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0101010100011)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==13'b0101010100100)) color_data = 12'b101000110011;
		if(({row_reg, col_reg}==13'b0101010100101)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==13'b0101010100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==13'b0101010100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0101010101000)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0101010101001)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0101010101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0101010101011)) color_data = 12'b010101010101;

		if(({row_reg, col_reg}>=13'b0101010101100) && ({row_reg, col_reg}<13'b0101011001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0101011001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b0101011001001) && ({row_reg, col_reg}<13'b0101011001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0101011001100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0101011001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=13'b0101011001110) && ({row_reg, col_reg}<13'b0101011010000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=13'b0101011010000) && ({row_reg, col_reg}<13'b0101011010010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0101011010010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0101011010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0101011010100) && ({row_reg, col_reg}<13'b0101011011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0101011011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==13'b0101011011101)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==13'b0101011011110)) color_data = 12'b101101010101;
		if(({row_reg, col_reg}>=13'b0101011011111) && ({row_reg, col_reg}<13'b0101011100001)) color_data = 12'b110001100110;
		if(({row_reg, col_reg}==13'b0101011100001)) color_data = 12'b101101000100;
		if(({row_reg, col_reg}==13'b0101011100010)) color_data = 12'b101000110011;
		if(({row_reg, col_reg}==13'b0101011100011)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==13'b0101011100100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==13'b0101011100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==13'b0101011100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0101011100111)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b0101011101000)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0101011101001)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b0101011101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0101011101011)) color_data = 12'b010001000100;

		if(({row_reg, col_reg}>=13'b0101011101100) && ({row_reg, col_reg}<13'b0101100001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0101100001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0101100001001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0101100001010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0101100001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0101100001100) && ({row_reg, col_reg}<13'b0101100001110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0101100001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0101100001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0101100010000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0101100010001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0101100010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0101100010011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0101100010100) && ({row_reg, col_reg}<13'b0101100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0101100011101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=13'b0101100011110) && ({row_reg, col_reg}<13'b0101100100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=13'b0101100100000) && ({row_reg, col_reg}<13'b0101100100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=13'b0101100100010) && ({row_reg, col_reg}<13'b0101100100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==13'b0101100100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==13'b0101100100101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0101100100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0101100100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0101100101000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0101100101001)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b0101100101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0101100101011)) color_data = 12'b001100110011;

		if(({row_reg, col_reg}>=13'b0101100101100) && ({row_reg, col_reg}<13'b0101101001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0101101001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0101101001001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0101101001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0101101001011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0101101001100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0101101001101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0101101001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0101101001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0101101010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0101101010001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0101101010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0101101010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=13'b0101101010100) && ({row_reg, col_reg}<13'b0101101100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0101101100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0101101100001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0101101100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0101101100011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0101101100100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0101101100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0101101100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0101101100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0101101101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0101101101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0101101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0101101101011)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=13'b0101101101100) && ({row_reg, col_reg}<13'b0101110001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0101110001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0101110001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0101110001010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0101110001011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=13'b0101110001100) && ({row_reg, col_reg}<13'b0101110001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0101110001110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0101110001111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0101110010000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0101110010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0101110010010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0101110010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0101110010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0101110010101) && ({row_reg, col_reg}<13'b0101110011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0101110011111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0101110100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0101110100001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0101110100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0101110100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0101110100100) && ({row_reg, col_reg}<13'b0101110100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0101110100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0101110100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0101110101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0101110101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0101110101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0101110101011)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=13'b0101110101100) && ({row_reg, col_reg}<13'b0101111001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0101111001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0101111001010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0101111001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0101111001100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0101111001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=13'b0101111001110) && ({row_reg, col_reg}<13'b0101111010000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0101111010000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0101111010001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0101111010010) && ({row_reg, col_reg}<13'b0101111010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0101111010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0101111010101) && ({row_reg, col_reg}<13'b0101111011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0101111011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0101111011111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0101111100000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0101111100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0101111100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0101111100011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=13'b0101111100100) && ({row_reg, col_reg}<13'b0101111100110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0101111100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0101111100111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0101111101000) && ({row_reg, col_reg}<13'b0101111101011)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=13'b0101111101011) && ({row_reg, col_reg}<13'b0110000001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0110000001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110000001010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0110000001011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0110000001100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0110000001101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0110000001110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0110000001111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0110000010000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0110000010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0110000010010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0110000010011) && ({row_reg, col_reg}<13'b0110000010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110000010101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0110000010110) && ({row_reg, col_reg}<13'b0110000011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0110000011110) && ({row_reg, col_reg}<13'b0110000100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110000100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0110000100010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0110000100011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=13'b0110000100100) && ({row_reg, col_reg}<13'b0110000100110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0110000100110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0110000100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0110000101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0110000101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110000101010)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=13'b0110000101011) && ({row_reg, col_reg}<13'b0110001001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0110001001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0110001001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110001001011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0110001001100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0110001001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0110001001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0110001001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0110001010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0110001010001) && ({row_reg, col_reg}<13'b0110001010011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0110001010011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0110001010100) && ({row_reg, col_reg}<13'b0110001010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b0110001010110) && ({row_reg, col_reg}<13'b0110001011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0110001011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110001011110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0110001011111) && ({row_reg, col_reg}<13'b0110001100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0110001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0110001100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0110001100011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0110001100100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0110001100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0110001100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0110001100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0110001101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110001101001)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=13'b0110001101010) && ({row_reg, col_reg}<13'b0110010001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0110010001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0110010001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110010001100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0110010001101) && ({row_reg, col_reg}<13'b0110010010001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0110010010001) && ({row_reg, col_reg}<13'b0110010010011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0110010010011) && ({row_reg, col_reg}<13'b0110010010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110010010101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0110010010110) && ({row_reg, col_reg}<13'b0110010011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0110010011101) && ({row_reg, col_reg}<13'b0110010011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0110010011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0110010100000) && ({row_reg, col_reg}<13'b0110010100010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0110010100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0110010100011) && ({row_reg, col_reg}<13'b0110010100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0110010100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0110010100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0110010100111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0110010101000)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=13'b0110010101001) && ({row_reg, col_reg}<13'b0110011001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0110011001010) && ({row_reg, col_reg}<13'b0110011001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b0110011001101) && ({row_reg, col_reg}<13'b0110011010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0110011010011) && ({row_reg, col_reg}<13'b0110011010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0110011010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0110011010110) && ({row_reg, col_reg}<13'b0110011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0110011011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110011011110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0110011011111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0110011100000) && ({row_reg, col_reg}<13'b0110011100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110011100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0110011100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0110011100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0110011100101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0110011100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0110011100111)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=13'b0110011101000) && ({row_reg, col_reg}<13'b0110100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0110100001011) && ({row_reg, col_reg}<13'b0110100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b0110100001101) && ({row_reg, col_reg}<13'b0110100001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110100001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0110100010000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0110100010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0110100010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0110100010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0110100010100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0110100010101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0110100010110) && ({row_reg, col_reg}<13'b0110100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0110100011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110100011110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0110100011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0110100100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0110100100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0110100100010) && ({row_reg, col_reg}<13'b0110100100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110100100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0110100100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110100100110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=13'b0110100100111) && ({row_reg, col_reg}<13'b0110101001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0110101001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0110101001110) && ({row_reg, col_reg}<13'b0110101010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0110101010011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0110101010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0110101010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0110101010110) && ({row_reg, col_reg}<13'b0110101011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0110101011101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0110101011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110101011111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0110101100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0110101100001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0110101100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0110101100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0110101100100) && ({row_reg, col_reg}<13'b0110101100110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=13'b0110101100110) && ({row_reg, col_reg}<13'b0110110001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0110110001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0110110001101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0110110001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0110110001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0110110010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0110110010001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0110110010010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0110110010011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0110110010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0110110010101) && ({row_reg, col_reg}<13'b0110110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0110110011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0110110011110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0110110011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110110100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0110110100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0110110100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0110110100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0110110100100)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=13'b0110110100101) && ({row_reg, col_reg}<13'b0110111001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0110111001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0110111001110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0110111001111) && ({row_reg, col_reg}<13'b0110111010010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0110111010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110111010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0110111010100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0110111010101) && ({row_reg, col_reg}<13'b0110111011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0110111011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110111011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0110111011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0110111100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110111100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0110111100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0110111100011)) color_data = 12'b010001000100;

		if(({row_reg, col_reg}>=13'b0110111100100) && ({row_reg, col_reg}<13'b0111000001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0111000001101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0111000001110) && ({row_reg, col_reg}<13'b0111000010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111000010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0111000010011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0111000010100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0111000010101) && ({row_reg, col_reg}<13'b0111000011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0111000011101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0111000011110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0111000011111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0111000100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0111000100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0111000100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111000100011)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=13'b0111000100100) && ({row_reg, col_reg}<13'b0111001001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0111001001101) && ({row_reg, col_reg}<13'b0111001001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0111001001111) && ({row_reg, col_reg}<13'b0111001010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0111001010001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0111001010010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0111001010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b0111001010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b0111001010101) && ({row_reg, col_reg}<13'b0111001011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0111001011101) && ({row_reg, col_reg}<13'b0111001011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111001011111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0111001100000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0111001100001) && ({row_reg, col_reg}<13'b0111001100011)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=13'b0111001100011) && ({row_reg, col_reg}<13'b0111010001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0111010001101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0111010001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0111010001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0111010010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111010010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0111010010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0111010010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0111010010100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0111010010101) && ({row_reg, col_reg}<13'b0111010011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0111010011100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0111010011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0111010011110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0111010011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111010100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0111010100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0111010100010) && ({row_reg, col_reg}<13'b0111010100100)) color_data = 12'b001100110011;

		if(({row_reg, col_reg}>=13'b0111010100100) && ({row_reg, col_reg}<13'b0111011001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0111011001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111011001110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0111011001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0111011010000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0111011010001) && ({row_reg, col_reg}<13'b0111011010011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0111011010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0111011010100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0111011010101) && ({row_reg, col_reg}<13'b0111011011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0111011011011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0111011011100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0111011011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0111011011110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0111011011111) && ({row_reg, col_reg}<13'b0111011100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111011100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0111011100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111011100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0111011100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0111011100101)) color_data = 12'b010101010101;

		if(({row_reg, col_reg}>=13'b0111011100110) && ({row_reg, col_reg}<13'b0111100001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0111100001100) && ({row_reg, col_reg}<13'b0111100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b0111100010001) && ({row_reg, col_reg}<13'b0111100010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0111100010101) && ({row_reg, col_reg}<13'b0111100011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0111100011011) && ({row_reg, col_reg}<13'b0111100011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0111100011101) && ({row_reg, col_reg}<13'b0111100011111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0111100011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0111100100000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0111100100001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0111100100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111100100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0111100100100) && ({row_reg, col_reg}<13'b0111100100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0111100100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0111100100111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0111100101000)) color_data = 12'b010101010101;

		if(({row_reg, col_reg}>=13'b0111100101001) && ({row_reg, col_reg}<13'b0111101001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0111101001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111101001100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0111101001101) && ({row_reg, col_reg}<13'b0111101001111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0111101001111) && ({row_reg, col_reg}<13'b0111101010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111101010001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0111101010010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0111101010011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0111101010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0111101010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0111101010110) && ({row_reg, col_reg}<13'b0111101011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0111101011010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0111101011011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0111101011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=13'b0111101011101) && ({row_reg, col_reg}<13'b0111101011111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0111101011111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0111101100000) && ({row_reg, col_reg}<13'b0111101100010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0111101100010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0111101100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0111101100100) && ({row_reg, col_reg}<13'b0111101100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111101100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0111101100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0111101101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0111101101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0111101101010)) color_data = 12'b001100110011;

		if(({row_reg, col_reg}>=13'b0111101101011) && ({row_reg, col_reg}<13'b0111110001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0111110001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0111110001011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0111110001100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0111110001101) && ({row_reg, col_reg}<13'b0111110001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0111110001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0111110010000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0111110010001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0111110010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0111110010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0111110010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0111110010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0111110010110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0111110010111) && ({row_reg, col_reg}<13'b0111110011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0111110011001)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0111110011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111110011011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0111110011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0111110011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0111110011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0111110011111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0111110100000)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b0111110100001)) color_data = 12'b110010010010;
		if(({row_reg, col_reg}==13'b0111110100010)) color_data = 12'b110110110100;
		if(({row_reg, col_reg}>=13'b0111110100011) && ({row_reg, col_reg}<13'b0111110100101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0111110100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0111110100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111110100111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0111110101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0111110101001)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0111110101010)) color_data = 12'b110010010010;
		if(({row_reg, col_reg}>=13'b0111110101011) && ({row_reg, col_reg}<13'b0111110101101)) color_data = 12'b111011010101;

		if(({row_reg, col_reg}>=13'b0111110101101) && ({row_reg, col_reg}<13'b0111111001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0111111001001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=13'b0111111001010) && ({row_reg, col_reg}<13'b0111111001100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0111111001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0111111001101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0111111001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111111001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0111111010000) && ({row_reg, col_reg}<13'b0111111010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111111010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0111111010100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b0111111010101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==13'b0111111010110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b0111111010111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0111111011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0111111011001)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0111111011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0111111011011) && ({row_reg, col_reg}<13'b0111111011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0111111011101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0111111011110) && ({row_reg, col_reg}<13'b0111111100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111111100000)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0111111100001)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0111111100010)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==13'b0111111100011)) color_data = 12'b110110110100;
		if(({row_reg, col_reg}>=13'b0111111100100) && ({row_reg, col_reg}<13'b0111111100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0111111100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b0111111100111) && ({row_reg, col_reg}<13'b0111111101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111111101001)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b0111111101010)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b0111111101011)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b0111111101100)) color_data = 12'b110110110100;
		if(({row_reg, col_reg}==13'b0111111101101)) color_data = 12'b110010010010;

		if(({row_reg, col_reg}>=13'b0111111101110) && ({row_reg, col_reg}<13'b1000000001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1000000001000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1000000001001) && ({row_reg, col_reg}<13'b1000000001011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1000000001011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b1000000001100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==13'b1000000001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b1000000001110) && ({row_reg, col_reg}<13'b1000000010001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1000000010001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1000000010010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b1000000010011) && ({row_reg, col_reg}<13'b1000000010101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b1000000010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b1000000010110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b1000000010111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1000000011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1000000011001)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}>=13'b1000000011010) && ({row_reg, col_reg}<13'b1000000011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b1000000011100) && ({row_reg, col_reg}<13'b1000000100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b1000000100000)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b1000000100001)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b1000000100010)) color_data = 12'b110010010010;
		if(({row_reg, col_reg}==13'b1000000100011)) color_data = 12'b110110110100;
		if(({row_reg, col_reg}==13'b1000000100100)) color_data = 12'b000100110000;
		if(({row_reg, col_reg}>=13'b1000000100101) && ({row_reg, col_reg}<13'b1000000101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1000000101000) && ({row_reg, col_reg}<13'b1000000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1000000101010)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}>=13'b1000000101011) && ({row_reg, col_reg}<13'b1000000101101)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b1000000101101)) color_data = 12'b010110100100;

		if(({row_reg, col_reg}>=13'b1000000101110) && ({row_reg, col_reg}<13'b1000001001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1000001001000)) color_data = 12'b110010010010;
		if(({row_reg, col_reg}==13'b1000001001001)) color_data = 12'b110110110100;
		if(({row_reg, col_reg}==13'b1000001001010)) color_data = 12'b110010010010;
		if(({row_reg, col_reg}==13'b1000001001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1000001001100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b1000001001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b1000001001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b1000001001111) && ({row_reg, col_reg}<13'b1000001010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1000001010001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1000001010010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b1000001010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b1000001010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1000001010101)) color_data = 12'b110010010010;
		if(({row_reg, col_reg}==13'b1000001010110)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==13'b1000001010111)) color_data = 12'b110010010010;
		if(({row_reg, col_reg}>=13'b1000001011000) && ({row_reg, col_reg}<13'b1000001100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1000001100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b1000001100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==13'b1000001100010)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b1000001100011)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}>=13'b1000001100100) && ({row_reg, col_reg}<13'b1000001101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1000001101101)) color_data = 12'b010010010011;

		if(({row_reg, col_reg}>=13'b1000001101110) && ({row_reg, col_reg}<13'b1000010000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1000010000111)) color_data = 12'b110010010010;
		if(({row_reg, col_reg}==13'b1000010001000)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==13'b1000010001001)) color_data = 12'b110010010010;
		if(({row_reg, col_reg}==13'b1000010001010)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b1000010001011)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b1000010001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1000010001101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1000010001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1000010001111) && ({row_reg, col_reg}<13'b1000010010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b1000010010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1000010010010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1000010010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1000010010100)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b1000010010101)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b1000010010110)) color_data = 12'b110110110100;
		if(({row_reg, col_reg}==13'b1000010010111)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==13'b1000010011000)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}>=13'b1000010011001) && ({row_reg, col_reg}<13'b1000010100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1000010100011)) color_data = 12'b010010010011;

		if(({row_reg, col_reg}>=13'b1000010100100) && ({row_reg, col_reg}<13'b1000011000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1000011000111)) color_data = 12'b110110110100;
		if(({row_reg, col_reg}==13'b1000011001000)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}>=13'b1000011001001) && ({row_reg, col_reg}<13'b1000011001011)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b1000011001011)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b1000011001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1000011001101) && ({row_reg, col_reg}<13'b1000011001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1000011001111) && ({row_reg, col_reg}<13'b1000011010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b1000011010010) && ({row_reg, col_reg}<13'b1000011010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b1000011010100)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==13'b1000011010101)) color_data = 12'b001110000010;
		if(({row_reg, col_reg}==13'b1000011010110)) color_data = 12'b010010010011;
		if(({row_reg, col_reg}==13'b1000011010111)) color_data = 12'b010110100100;
		if(({row_reg, col_reg}==13'b1000011011000)) color_data = 12'b110010010010;

		if(({row_reg, col_reg}>=13'b1000011011001) && ({row_reg, col_reg}<13'b1000100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1000100000111)) color_data = 12'b110010010010;
		if(({row_reg, col_reg}>=13'b1000100001000) && ({row_reg, col_reg}<13'b1000100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1000100011000)) color_data = 12'b110010010010;

		if(({row_reg, col_reg}>=13'b1000100011001) && ({row_reg, col_reg}<=13'b1000100110001)) color_data = 12'b000000000000;
	end
endmodule