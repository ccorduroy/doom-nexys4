module bgr_rom
	(
		input wire clk,
		input wire [7:0] row,
		input wire [7:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [7:0] row_reg;
	reg [7:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin
		if(({row_reg, col_reg}==16'b0000000000000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000000000000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000000000000010) && ({row_reg, col_reg}<16'b0000000000000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000000000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000000000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000000000001000) && ({row_reg, col_reg}<16'b0000000000001010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000000000001010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000000001011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000000000001100) && ({row_reg, col_reg}<16'b0000000000001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000000001110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000000000001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000000010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000000010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000000000010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000000000010011) && ({row_reg, col_reg}<16'b0000000000010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000000010101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000000000010110) && ({row_reg, col_reg}<16'b0000000000011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000000000011011) && ({row_reg, col_reg}<16'b0000000000011101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000000000011101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000000000011110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000000000011111) && ({row_reg, col_reg}<16'b0000000000100111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000000000100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000000101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000000101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000000000101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000000101011) && ({row_reg, col_reg}<16'b0000000000101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000000101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000000101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000000101111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000000000110000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000000000110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000000000110010) && ({row_reg, col_reg}<16'b0000000000110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000000000110100) && ({row_reg, col_reg}<16'b0000000000110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000000110110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000000000110111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000000000111000) && ({row_reg, col_reg}<16'b0000000000111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000000111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000000000111011) && ({row_reg, col_reg}<16'b0000000000111101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000000000111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000000111110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000000000111111) && ({row_reg, col_reg}<16'b0000000001000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000000001000001) && ({row_reg, col_reg}<16'b0000000001000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000000001000101) && ({row_reg, col_reg}<16'b0000000001000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000001000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000000001001000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000000001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000000001001010) && ({row_reg, col_reg}<16'b0000000001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000001001100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000000001001101) && ({row_reg, col_reg}<16'b0000000001010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000001010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000000001010001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0000000001010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000000001010011) && ({row_reg, col_reg}<16'b0000000001010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000001010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000001011000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0000000001011001) && ({row_reg, col_reg}<16'b0000000001011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000000001011101) && ({row_reg, col_reg}<16'b0000000001100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000000001100000) && ({row_reg, col_reg}<16'b0000000001100010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000000001100010) && ({row_reg, col_reg}<16'b0000000001100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000000001100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000000001100110) && ({row_reg, col_reg}<16'b0000000001101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000000001101000) && ({row_reg, col_reg}<16'b0000000001101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000000001101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000001101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000000001101110) && ({row_reg, col_reg}<16'b0000000001110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000000001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000001110001) && ({row_reg, col_reg}<16'b0000000001110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000000001110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000000001110100) && ({row_reg, col_reg}<16'b0000000001110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000001110110) && ({row_reg, col_reg}<16'b0000000001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000001111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000000001111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000000001111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000000001111011) && ({row_reg, col_reg}<16'b0000000010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000010000011) && ({row_reg, col_reg}<16'b0000000010100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000000010100010) && ({row_reg, col_reg}<16'b0000000010100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000000010100110) && ({row_reg, col_reg}<16'b0000000010101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000000010101011) && ({row_reg, col_reg}<16'b0000000010101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000000010101101) && ({row_reg, col_reg}<16'b0000000010110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000010110010) && ({row_reg, col_reg}<16'b0000000010110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000000010110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000000010110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000000010110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000010110111) && ({row_reg, col_reg}<16'b0000000011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000000011000001) && ({row_reg, col_reg}<16'b0000000011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000011001110) && ({row_reg, col_reg}<16'b0000000011010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000000011010000) && ({row_reg, col_reg}<16'b0000000011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000011011111) && ({row_reg, col_reg}<16'b0000000011100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000000011100011) && ({row_reg, col_reg}<16'b0000000011100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000011100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000011100110) && ({row_reg, col_reg}<16'b0000000011101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000000011101100) && ({row_reg, col_reg}<16'b0000000011101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000011101110) && ({row_reg, col_reg}<16'b0000000011110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000000011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000011110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000011110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000011110100) && ({row_reg, col_reg}<16'b0000000011110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000011110111) && ({row_reg, col_reg}<16'b0000000011111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000011111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000011111010) && ({row_reg, col_reg}<16'b0000000011111110)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0000000011111110) && ({row_reg, col_reg}<16'b0000000100000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000100000000) && ({row_reg, col_reg}<16'b0000000100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000100000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000000100000011) && ({row_reg, col_reg}<16'b0000000100000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000100000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000000100000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000100000111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000000100001000) && ({row_reg, col_reg}<16'b0000000100001010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000000100001010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000000100001011) && ({row_reg, col_reg}<16'b0000000100001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000100001110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000000100001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000100010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000100010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000000100010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000000100010011) && ({row_reg, col_reg}<16'b0000000100010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000000100010101) && ({row_reg, col_reg}<16'b0000000100010111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000100010111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0000000100011000) && ({row_reg, col_reg}<16'b0000000100100100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000000100100100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000000100100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000100100110)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000000100100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000100101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000100101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000000100101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000100101011) && ({row_reg, col_reg}<16'b0000000100101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000100101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000100101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000000100101111) && ({row_reg, col_reg}<16'b0000000100110001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000000100110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000000100110010) && ({row_reg, col_reg}<16'b0000000100110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000000100110100) && ({row_reg, col_reg}<16'b0000000100110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000100110111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000000100111000) && ({row_reg, col_reg}<16'b0000000100111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000100111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000000100111011) && ({row_reg, col_reg}<16'b0000000100111101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000000100111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000100111110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000000100111111) && ({row_reg, col_reg}<16'b0000000101000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000000101000001) && ({row_reg, col_reg}<16'b0000000101000110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000000101000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000000101000111) && ({row_reg, col_reg}<16'b0000000101001001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000000101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000000101001010) && ({row_reg, col_reg}<16'b0000000101001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000000101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000101001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000101001110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000000101001111) && ({row_reg, col_reg}<16'b0000000101010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000000101010011) && ({row_reg, col_reg}<16'b0000000101010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000000101010110) && ({row_reg, col_reg}<16'b0000000101011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000000101011001) && ({row_reg, col_reg}<16'b0000000101100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000101100010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000000101100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0000000101100100) && ({row_reg, col_reg}<16'b0000000101100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000000101100110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000000101100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000000101101000) && ({row_reg, col_reg}<16'b0000000101101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000000101101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000000101101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000101101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000101101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000000101101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000000101110000) && ({row_reg, col_reg}<16'b0000000101110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000101110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000000101110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000000101110100) && ({row_reg, col_reg}<16'b0000000101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000101110110) && ({row_reg, col_reg}<16'b0000000101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000101111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000000101111001) && ({row_reg, col_reg}<16'b0000000101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000101111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000101111101) && ({row_reg, col_reg}<16'b0000000110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000110000011) && ({row_reg, col_reg}<16'b0000000110100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000000110100011) && ({row_reg, col_reg}<16'b0000000110100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000110100110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000110100111) && ({row_reg, col_reg}<16'b0000000110101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000000110101011) && ({row_reg, col_reg}<16'b0000000110101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000000110101101) && ({row_reg, col_reg}<16'b0000000110110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000110110011) && ({row_reg, col_reg}<16'b0000000110110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000000110110111) && ({row_reg, col_reg}<16'b0000000110111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000110111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000110111010) && ({row_reg, col_reg}<16'b0000000110111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000110111111) && ({row_reg, col_reg}<16'b0000000111000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000000111000001) && ({row_reg, col_reg}<16'b0000000111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000111001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000000111001010) && ({row_reg, col_reg}<16'b0000000111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000111001110) && ({row_reg, col_reg}<16'b0000000111010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000000111010000) && ({row_reg, col_reg}<16'b0000000111010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000111010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000000111010111) && ({row_reg, col_reg}<16'b0000000111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000111011111) && ({row_reg, col_reg}<16'b0000000111100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000000111100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000111100100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000111100101) && ({row_reg, col_reg}<16'b0000000111100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000000111100111) && ({row_reg, col_reg}<16'b0000000111101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000000111101011) && ({row_reg, col_reg}<16'b0000000111101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000000111101101) && ({row_reg, col_reg}<16'b0000000111110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000000111110001) && ({row_reg, col_reg}<16'b0000000111111001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0000000111111001) && ({row_reg, col_reg}<16'b0000001000000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001000000000) && ({row_reg, col_reg}<16'b0000001000000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000001000000011) && ({row_reg, col_reg}<16'b0000001000000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001000000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000001000000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001000000111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000001000001000) && ({row_reg, col_reg}<16'b0000001000001010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000001000001010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001000001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001000001100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000001000001101) && ({row_reg, col_reg}<16'b0000001000010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001000010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001000010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001000010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000001000010011) && ({row_reg, col_reg}<16'b0000001000010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000001000010101) && ({row_reg, col_reg}<16'b0000001000011000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000001000011000) && ({row_reg, col_reg}<16'b0000001000100100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000001000100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001000100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000001000100110) && ({row_reg, col_reg}<16'b0000001000101000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001000101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001000101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000001000101010) && ({row_reg, col_reg}<16'b0000001000101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001000101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001000101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000001000101111) && ({row_reg, col_reg}<16'b0000001000110001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000001000110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001000110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001000110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000001000110100) && ({row_reg, col_reg}<16'b0000001000110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001000110111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000001000111000) && ({row_reg, col_reg}<16'b0000001000111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001000111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000001000111011) && ({row_reg, col_reg}<16'b0000001000111101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000001000111101) && ({row_reg, col_reg}<16'b0000001001000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000001001000000) && ({row_reg, col_reg}<16'b0000001001000100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000001001000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001001000101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000001001000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000001001000111) && ({row_reg, col_reg}<16'b0000001001001001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001001001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001001001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000001001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001001001101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000001001001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000001001001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000001001010000) && ({row_reg, col_reg}<16'b0000001001010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000001001010011) && ({row_reg, col_reg}<16'b0000001001010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001001010101)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0000001001010110) && ({row_reg, col_reg}<16'b0000001001011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000001001011001) && ({row_reg, col_reg}<16'b0000001001011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001001011100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000001001011101) && ({row_reg, col_reg}<16'b0000001001100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001001100001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000001001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000001001100011) && ({row_reg, col_reg}<16'b0000001001100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000001001100111) && ({row_reg, col_reg}<16'b0000001001101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000001001101001) && ({row_reg, col_reg}<16'b0000001001101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000001001101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001001101100) && ({row_reg, col_reg}<16'b0000001001101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001001101110) && ({row_reg, col_reg}<16'b0000001001110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000001001110000) && ({row_reg, col_reg}<16'b0000001001110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001001110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000001001110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000001001110100) && ({row_reg, col_reg}<16'b0000001001110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001001110110) && ({row_reg, col_reg}<16'b0000001001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001001111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000001001111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001001111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000001001111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000001001111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000001001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000001001111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000001010000000) && ({row_reg, col_reg}<16'b0000001010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001010000011) && ({row_reg, col_reg}<16'b0000001010100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000001010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001010100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000001010100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001010100110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001010100111) && ({row_reg, col_reg}<16'b0000001010101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000001010101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001010101011) && ({row_reg, col_reg}<16'b0000001010101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000001010101101) && ({row_reg, col_reg}<16'b0000001010110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001010110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001010110010) && ({row_reg, col_reg}<16'b0000001010110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001010110100) && ({row_reg, col_reg}<16'b0000001010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000001010110110) && ({row_reg, col_reg}<16'b0000001010111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000001011000000) && ({row_reg, col_reg}<16'b0000001011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001011001000) && ({row_reg, col_reg}<16'b0000001011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000001011001011) && ({row_reg, col_reg}<16'b0000001011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001011001110) && ({row_reg, col_reg}<16'b0000001011010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000001011010000) && ({row_reg, col_reg}<16'b0000001011100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001011100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000001011100110) && ({row_reg, col_reg}<16'b0000001011101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001011101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000001011101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000001011101011) && ({row_reg, col_reg}<16'b0000001011101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001011101101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0000001011101110) && ({row_reg, col_reg}<16'b0000001011110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000001011110000) && ({row_reg, col_reg}<16'b0000001011110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001011110100) && ({row_reg, col_reg}<16'b0000001011110111)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0000001011110111) && ({row_reg, col_reg}<16'b0000001100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000001100000001) && ({row_reg, col_reg}<16'b0000001100000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000001100000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000001100000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001100000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001100000110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000001100000111)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000001100001000)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==16'b0000001100001001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000001100001010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001100001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001100001100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000001100001101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000001100001110) && ({row_reg, col_reg}<16'b0000001100010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001100010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001100010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001100010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000001100010011) && ({row_reg, col_reg}<16'b0000001100010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000001100010101) && ({row_reg, col_reg}<16'b0000001100010111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000001100010111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000001100011000) && ({row_reg, col_reg}<16'b0000001100100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001100100011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000001100100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000001100100101) && ({row_reg, col_reg}<16'b0000001100101000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000001100101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001100101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001100101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000001100101011) && ({row_reg, col_reg}<16'b0000001100101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001100101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001100101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000001100101111) && ({row_reg, col_reg}<16'b0000001100110001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001100110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001100110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001100110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000001100110100) && ({row_reg, col_reg}<16'b0000001100110110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000001100110110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000001100110111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000001100111000) && ({row_reg, col_reg}<16'b0000001100111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001100111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000001100111011) && ({row_reg, col_reg}<16'b0000001100111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000001100111101) && ({row_reg, col_reg}<16'b0000001100111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000001100111111) && ({row_reg, col_reg}<16'b0000001101000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000001101000011) && ({row_reg, col_reg}<16'b0000001101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001101000110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0000001101000111)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0000001101001000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001101001001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000001101001010) && ({row_reg, col_reg}<16'b0000001101001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001101001101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000001101001110) && ({row_reg, col_reg}<16'b0000001101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001101010000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0000001101010001) && ({row_reg, col_reg}<16'b0000001101010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000001101010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001101010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000001101010101) && ({row_reg, col_reg}<16'b0000001101100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001101100000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000001101100001) && ({row_reg, col_reg}<16'b0000001101100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000001101100011) && ({row_reg, col_reg}<16'b0000001101100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001101100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000001101100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001101100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000001101101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001101101001) && ({row_reg, col_reg}<16'b0000001101101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001101101100) && ({row_reg, col_reg}<16'b0000001101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001101101110) && ({row_reg, col_reg}<16'b0000001101110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000001101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001101110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001101110010) && ({row_reg, col_reg}<16'b0000001101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000001101110100) && ({row_reg, col_reg}<16'b0000001101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001101110110) && ({row_reg, col_reg}<16'b0000001101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001101111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000001101111001) && ({row_reg, col_reg}<16'b0000001101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000001101111011)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==16'b0000001101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000001101111101) && ({row_reg, col_reg}<16'b0000001110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001110000000) && ({row_reg, col_reg}<16'b0000001110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001110000011) && ({row_reg, col_reg}<16'b0000001110100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000001110100100) && ({row_reg, col_reg}<16'b0000001110100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001110100110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001110100111) && ({row_reg, col_reg}<16'b0000001110101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000001110101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001110101011) && ({row_reg, col_reg}<16'b0000001110101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000001110101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000001110101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000001110110000) && ({row_reg, col_reg}<16'b0000001110110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001110110011) && ({row_reg, col_reg}<16'b0000001110111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001110111011) && ({row_reg, col_reg}<16'b0000001110111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000001110111101) && ({row_reg, col_reg}<16'b0000001111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001111000111) && ({row_reg, col_reg}<16'b0000001111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000001111001011) && ({row_reg, col_reg}<16'b0000001111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001111001110) && ({row_reg, col_reg}<16'b0000001111010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000001111010001) && ({row_reg, col_reg}<16'b0000001111011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001111011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000001111011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001111011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000001111011101) && ({row_reg, col_reg}<16'b0000001111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001111011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000001111100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000001111100001) && ({row_reg, col_reg}<16'b0000001111100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001111100100) && ({row_reg, col_reg}<16'b0000001111100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000001111100110) && ({row_reg, col_reg}<16'b0000001111101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001111101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000001111101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000001111101100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0000001111101101) && ({row_reg, col_reg}<16'b0000001111110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000001111110000) && ({row_reg, col_reg}<16'b0000001111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001111110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001111110011) && ({row_reg, col_reg}<16'b0000001111110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000001111110110) && ({row_reg, col_reg}<16'b0000001111111000)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0000001111111000) && ({row_reg, col_reg}<16'b0000010000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000010000000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010000000010) && ({row_reg, col_reg}<16'b0000010000000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000010000000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010000000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010000000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010000000111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000010000001000) && ({row_reg, col_reg}<16'b0000010000001010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000010000001010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000010000001011) && ({row_reg, col_reg}<16'b0000010000001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010000001110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000010000001111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000010000010000) && ({row_reg, col_reg}<16'b0000010000010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010000010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000010000010011) && ({row_reg, col_reg}<16'b0000010000011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000010000011010) && ({row_reg, col_reg}<16'b0000010000011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000010000011100) && ({row_reg, col_reg}<16'b0000010000100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010000100000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000010000100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010000100010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000010000100011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000010000100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010000100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000010000100110) && ({row_reg, col_reg}<16'b0000010000101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010000101000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000010000101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010000101010) && ({row_reg, col_reg}<16'b0000010000101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000010000101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010000101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000010000101111) && ({row_reg, col_reg}<16'b0000010000110001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010000110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000010000110010) && ({row_reg, col_reg}<16'b0000010000110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000010000110100) && ({row_reg, col_reg}<16'b0000010000110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010000110110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0000010000110111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000010000111000) && ({row_reg, col_reg}<16'b0000010000111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010000111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000010000111011) && ({row_reg, col_reg}<16'b0000010000111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010000111101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000010000111110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000010000111111) && ({row_reg, col_reg}<16'b0000010001000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000010001000011) && ({row_reg, col_reg}<16'b0000010001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010001000101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000010001000110) && ({row_reg, col_reg}<16'b0000010001001001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0000010001001001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000010001001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000010001001011) && ({row_reg, col_reg}<16'b0000010001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010001010000) && ({row_reg, col_reg}<16'b0000010001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000010001010100) && ({row_reg, col_reg}<16'b0000010001011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010001011001) && ({row_reg, col_reg}<16'b0000010001011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010001011100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0000010001011101) && ({row_reg, col_reg}<16'b0000010001011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000010001011111) && ({row_reg, col_reg}<16'b0000010001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010001100010) && ({row_reg, col_reg}<16'b0000010001100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010001100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000010001101000) && ({row_reg, col_reg}<16'b0000010001101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010001101110) && ({row_reg, col_reg}<16'b0000010001110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000010001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010001110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010001110010) && ({row_reg, col_reg}<16'b0000010001110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000010001110100) && ({row_reg, col_reg}<16'b0000010001110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010001110110) && ({row_reg, col_reg}<16'b0000010001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010001111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000010001111001) && ({row_reg, col_reg}<16'b0000010001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010001111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010001111100) && ({row_reg, col_reg}<16'b0000010001111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000010001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010010000000) && ({row_reg, col_reg}<16'b0000010010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010010000011) && ({row_reg, col_reg}<16'b0000010010101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000010010101011) && ({row_reg, col_reg}<16'b0000010010101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000010010101110) && ({row_reg, col_reg}<16'b0000010010110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010010110100) && ({row_reg, col_reg}<16'b0000010010111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010010111011) && ({row_reg, col_reg}<16'b0000010010111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000010010111101) && ({row_reg, col_reg}<16'b0000010010111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010010111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010011000000) && ({row_reg, col_reg}<16'b0000010011000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010011000110) && ({row_reg, col_reg}<16'b0000010011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000010011001010) && ({row_reg, col_reg}<16'b0000010011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010011001110) && ({row_reg, col_reg}<16'b0000010011010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000010011010001) && ({row_reg, col_reg}<16'b0000010011010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010011010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010011010101) && ({row_reg, col_reg}<16'b0000010011011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010011011001) && ({row_reg, col_reg}<16'b0000010011011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000010011011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000010011100000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=16'b0000010011100001) && ({row_reg, col_reg}<16'b0000010011100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010011100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000010011100100) && ({row_reg, col_reg}<16'b0000010011100110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000010011100110) && ({row_reg, col_reg}<16'b0000010011101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000010011101001) && ({row_reg, col_reg}<16'b0000010011101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010011101011) && ({row_reg, col_reg}<16'b0000010011110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000010011110000) && ({row_reg, col_reg}<16'b0000010011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010011110010) && ({row_reg, col_reg}<16'b0000010011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000010011111000)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0000010011111001) && ({row_reg, col_reg}<16'b0000010100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000010100000001) && ({row_reg, col_reg}<16'b0000010100000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000010100000011) && ({row_reg, col_reg}<16'b0000010100000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010100000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010100000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010100000111)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0000010100001000) && ({row_reg, col_reg}<16'b0000010100001010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0000010100001010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000010100001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000010100001100) && ({row_reg, col_reg}<16'b0000010100010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010100010010) && ({row_reg, col_reg}<16'b0000010100010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000010100010100) && ({row_reg, col_reg}<16'b0000010100011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010100011001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000010100011010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010100011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000010100011100) && ({row_reg, col_reg}<16'b0000010100100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010100100000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000010100100001) && ({row_reg, col_reg}<16'b0000010100100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000010100100011) && ({row_reg, col_reg}<16'b0000010100100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000010100100101) && ({row_reg, col_reg}<16'b0000010100101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000010100101001) && ({row_reg, col_reg}<16'b0000010100101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010100101011) && ({row_reg, col_reg}<16'b0000010100101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000010100101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010100101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000010100101111) && ({row_reg, col_reg}<16'b0000010100110001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010100110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010100110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000010100110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000010100110100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0000010100110101) && ({row_reg, col_reg}<16'b0000010100110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000010100110111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000010100111000) && ({row_reg, col_reg}<16'b0000010100111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010100111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010100111011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000010100111100) && ({row_reg, col_reg}<16'b0000010100111110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010100111110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000010100111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010101000000) && ({row_reg, col_reg}<16'b0000010101000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000010101000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010101000100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000010101000101) && ({row_reg, col_reg}<16'b0000010101000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000010101000111) && ({row_reg, col_reg}<16'b0000010101001001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000010101001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0000010101001010) && ({row_reg, col_reg}<16'b0000010101001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000010101001101) && ({row_reg, col_reg}<16'b0000010101001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010101001111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0000010101010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000010101010001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0000010101010010) && ({row_reg, col_reg}<16'b0000010101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000010101010100) && ({row_reg, col_reg}<16'b0000010101011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010101011001) && ({row_reg, col_reg}<16'b0000010101011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000010101011011) && ({row_reg, col_reg}<16'b0000010101100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010101100001) && ({row_reg, col_reg}<16'b0000010101100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010101100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000010101100100) && ({row_reg, col_reg}<16'b0000010101100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010101100110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000010101100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000010101101000) && ({row_reg, col_reg}<16'b0000010101101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010101101101) && ({row_reg, col_reg}<16'b0000010101110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000010101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010101110001) && ({row_reg, col_reg}<16'b0000010101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000010101110100) && ({row_reg, col_reg}<16'b0000010101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010101110110) && ({row_reg, col_reg}<16'b0000010101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010101111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000010101111001) && ({row_reg, col_reg}<16'b0000010101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010101111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000010101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000010101111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000010101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000010101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010110000000) && ({row_reg, col_reg}<16'b0000010110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010110000011) && ({row_reg, col_reg}<16'b0000010110101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000010110101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010110101100) && ({row_reg, col_reg}<16'b0000010110101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000010110101110) && ({row_reg, col_reg}<16'b0000010110110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010110110011) && ({row_reg, col_reg}<16'b0000010110110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010110110110) && ({row_reg, col_reg}<16'b0000010110111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010110111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000010110111101) && ({row_reg, col_reg}<16'b0000010111000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010111000010) && ({row_reg, col_reg}<16'b0000010111000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000010111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010111000110) && ({row_reg, col_reg}<16'b0000010111001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000010111001000) && ({row_reg, col_reg}<16'b0000010111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010111001110) && ({row_reg, col_reg}<16'b0000010111010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000010111010000) && ({row_reg, col_reg}<16'b0000010111010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010111010011) && ({row_reg, col_reg}<16'b0000010111010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010111010101) && ({row_reg, col_reg}<16'b0000010111011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010111011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000010111011010)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=16'b0000010111011011) && ({row_reg, col_reg}<16'b0000010111100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000010111100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010111100011) && ({row_reg, col_reg}<16'b0000010111101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000010111101001) && ({row_reg, col_reg}<16'b0000010111101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010111101110) && ({row_reg, col_reg}<16'b0000010111110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000010111110000) && ({row_reg, col_reg}<16'b0000010111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010111110010) && ({row_reg, col_reg}<16'b0000010111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000010111111001)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0000010111111010) && ({row_reg, col_reg}<16'b0000011000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011000000000) && ({row_reg, col_reg}<16'b0000011000000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011000000010) && ({row_reg, col_reg}<16'b0000011000000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0000011000000100) && ({row_reg, col_reg}<16'b0000011000000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011000000110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0000011000000111) && ({row_reg, col_reg}<16'b0000011000001001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000011000001001) && ({row_reg, col_reg}<16'b0000011000001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0000011000001011) && ({row_reg, col_reg}<16'b0000011000001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000011000001101) && ({row_reg, col_reg}<16'b0000011000010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000011000010010) && ({row_reg, col_reg}<16'b0000011000010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000011000010101) && ({row_reg, col_reg}<16'b0000011000011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000011000011000) && ({row_reg, col_reg}<16'b0000011000011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011000011100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000011000011101) && ({row_reg, col_reg}<16'b0000011000011111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000011000011111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000011000100000) && ({row_reg, col_reg}<16'b0000011000100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011000100101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0000011000100110) && ({row_reg, col_reg}<16'b0000011000101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011000101000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000011000101001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000011000101010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000011000101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011000101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000011000101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011000101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000011000101111) && ({row_reg, col_reg}<16'b0000011000110001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011000110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011000110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000011000110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000011000110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0000011000110101) && ({row_reg, col_reg}<16'b0000011000110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000011000110111) && ({row_reg, col_reg}<16'b0000011000111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011000111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011000111011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000011000111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000011000111101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000011000111110) && ({row_reg, col_reg}<16'b0000011001000000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000011001000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000011001000001) && ({row_reg, col_reg}<16'b0000011001000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000011001000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011001000100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000011001000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011001000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000011001001000) && ({row_reg, col_reg}<16'b0000011001001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000011001001010)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b0000011001001011) && ({row_reg, col_reg}<16'b0000011001001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000011001001101)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}==16'b0000011001001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011001001111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0000011001010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000011001010001)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0000011001010010)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0000011001010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000011001010100) && ({row_reg, col_reg}<16'b0000011001010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011001010111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000011001011000) && ({row_reg, col_reg}<16'b0000011001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000011001100010) && ({row_reg, col_reg}<16'b0000011001100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000011001100110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0000011001100111) && ({row_reg, col_reg}<16'b0000011001101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000011001101001) && ({row_reg, col_reg}<16'b0000011001101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011001101011) && ({row_reg, col_reg}<16'b0000011001101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011001101101) && ({row_reg, col_reg}<16'b0000011001110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000011001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011001110001) && ({row_reg, col_reg}<16'b0000011001110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000011001110100) && ({row_reg, col_reg}<16'b0000011001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011001111000) && ({row_reg, col_reg}<16'b0000011001111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000011001111010) && ({row_reg, col_reg}<16'b0000011001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011001111100) && ({row_reg, col_reg}<16'b0000011001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000011001111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000011010000000) && ({row_reg, col_reg}<16'b0000011010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011010000011) && ({row_reg, col_reg}<16'b0000011010101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000011010101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011010101101) && ({row_reg, col_reg}<16'b0000011010110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000011010110100) && ({row_reg, col_reg}<16'b0000011010110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011010110110) && ({row_reg, col_reg}<16'b0000011011000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011011000110) && ({row_reg, col_reg}<16'b0000011011001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011011001000) && ({row_reg, col_reg}<16'b0000011011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011011001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011011001011) && ({row_reg, col_reg}<16'b0000011011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011011001110) && ({row_reg, col_reg}<16'b0000011011010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000011011010000) && ({row_reg, col_reg}<16'b0000011011010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011011010011) && ({row_reg, col_reg}<16'b0000011011010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011011010101) && ({row_reg, col_reg}<16'b0000011011010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011011010111) && ({row_reg, col_reg}<16'b0000011011011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011011011100) && ({row_reg, col_reg}<16'b0000011011100010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000011011100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011011100011) && ({row_reg, col_reg}<16'b0000011011110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000011011110000) && ({row_reg, col_reg}<16'b0000011011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011011110010) && ({row_reg, col_reg}<16'b0000011011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000011011111001) && ({row_reg, col_reg}<16'b0000011011111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0000011011111011) && ({row_reg, col_reg}<16'b0000011100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011100000000) && ({row_reg, col_reg}<16'b0000011100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011100000010) && ({row_reg, col_reg}<16'b0000011100000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0000011100000100) && ({row_reg, col_reg}<16'b0000011100000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011100000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000011100001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000011100001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011100001010) && ({row_reg, col_reg}<16'b0000011100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000011100001100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000011100001101) && ({row_reg, col_reg}<16'b0000011100001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000011100001111) && ({row_reg, col_reg}<16'b0000011100010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000011100010001) && ({row_reg, col_reg}<16'b0000011100010011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0000011100010011) && ({row_reg, col_reg}<16'b0000011100010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000011100010101) && ({row_reg, col_reg}<16'b0000011100011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011100011000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000011100011001) && ({row_reg, col_reg}<16'b0000011100100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000011100100001) && ({row_reg, col_reg}<16'b0000011100100100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000011100100100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0000011100100101) && ({row_reg, col_reg}<16'b0000011100101000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0000011100101000) && ({row_reg, col_reg}<16'b0000011100101010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000011100101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011100101011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000011100101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011100101101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000011100101110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000011100101111)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000011100110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011100110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000011100110010) && ({row_reg, col_reg}<16'b0000011100110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000011100110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000011100110101) && ({row_reg, col_reg}<16'b0000011100110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000011100110111) && ({row_reg, col_reg}<16'b0000011100111001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011100111001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000011100111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000011100111011) && ({row_reg, col_reg}<16'b0000011100111101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000011100111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011100111110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000011100111111) && ({row_reg, col_reg}<16'b0000011101000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000011101000001) && ({row_reg, col_reg}<16'b0000011101000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000011101000011) && ({row_reg, col_reg}<16'b0000011101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011101000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000011101000111) && ({row_reg, col_reg}<16'b0000011101001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000011101001001)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==16'b0000011101001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000011101001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000011101001100) && ({row_reg, col_reg}<16'b0000011101001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000011101001111) && ({row_reg, col_reg}<16'b0000011101010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000011101010001)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0000011101010010)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0000011101010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000011101010100) && ({row_reg, col_reg}<16'b0000011101010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000011101010111) && ({row_reg, col_reg}<16'b0000011101011010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000011101011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000011101011011) && ({row_reg, col_reg}<16'b0000011101011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000011101011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011101011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000011101011111) && ({row_reg, col_reg}<16'b0000011101100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011101100010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0000011101100011) && ({row_reg, col_reg}<16'b0000011101100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000011101100111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0000011101101000) && ({row_reg, col_reg}<16'b0000011101101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000011101101010) && ({row_reg, col_reg}<16'b0000011101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011101101111) && ({row_reg, col_reg}<16'b0000011101110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011101110001) && ({row_reg, col_reg}<16'b0000011101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000011101110100) && ({row_reg, col_reg}<16'b0000011101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011101110110) && ({row_reg, col_reg}<16'b0000011101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011101111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000011101111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000011101111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011101111011) && ({row_reg, col_reg}<16'b0000011101111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000011101111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000011110000000) && ({row_reg, col_reg}<16'b0000011110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011110000011) && ({row_reg, col_reg}<16'b0000011110101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000011110101011) && ({row_reg, col_reg}<16'b0000011110101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011110101101) && ({row_reg, col_reg}<16'b0000011110110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011110110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011110110011) && ({row_reg, col_reg}<16'b0000011110110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000011110110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011110110110) && ({row_reg, col_reg}<16'b0000011110111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011110111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011111000000) && ({row_reg, col_reg}<16'b0000011111000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011111000110) && ({row_reg, col_reg}<16'b0000011111001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011111001000) && ({row_reg, col_reg}<16'b0000011111010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011111010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000011111010001) && ({row_reg, col_reg}<16'b0000011111010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011111010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011111010101) && ({row_reg, col_reg}<16'b0000011111010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011111010111) && ({row_reg, col_reg}<16'b0000011111011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000011111011011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000011111011100) && ({row_reg, col_reg}<16'b0000011111011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000011111011111) && ({row_reg, col_reg}<16'b0000011111101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000011111101011) && ({row_reg, col_reg}<16'b0000011111101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000011111101101) && ({row_reg, col_reg}<16'b0000011111110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000011111110000) && ({row_reg, col_reg}<16'b0000011111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011111110010) && ({row_reg, col_reg}<16'b0000011111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000011111111001) && ({row_reg, col_reg}<16'b0000011111111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0000011111111011) && ({row_reg, col_reg}<16'b0000100000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000100000000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000100000000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100000000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0000100000000100) && ({row_reg, col_reg}<16'b0000100000000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100000000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100000001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100000001001) && ({row_reg, col_reg}<16'b0000100000001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000100000001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000100000001100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000100000001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100000001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000100000001111) && ({row_reg, col_reg}<16'b0000100000010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000100000010001)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0000100000010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0000100000010011) && ({row_reg, col_reg}<16'b0000100000010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000100000010101) && ({row_reg, col_reg}<16'b0000100000011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100000011001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000100000011010) && ({row_reg, col_reg}<16'b0000100000100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100000100001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000100000100010)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0000100000100011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000100000100100)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0000100000100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100000100110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0000100000100111)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0000100000101000)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0000100000101001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000100000101010)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0000100000101011) && ({row_reg, col_reg}<16'b0000100000101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100000101110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100000101111)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000100000110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100000110001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000100000110010) && ({row_reg, col_reg}<16'b0000100000110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000100000110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100000110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100000110110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000100000110111) && ({row_reg, col_reg}<16'b0000100000111001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100000111001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000100000111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100000111011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000100000111100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000100000111101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100000111110)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000100000111111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000100001000000)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0000100001000001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0000100001000010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000100001000011) && ({row_reg, col_reg}<16'b0000100001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100001000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000100001000111) && ({row_reg, col_reg}<16'b0000100001001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000100001001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000100001001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000100001001100) && ({row_reg, col_reg}<16'b0000100001001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000100001001111) && ({row_reg, col_reg}<16'b0000100001010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000100001010001)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}>=16'b0000100001010010) && ({row_reg, col_reg}<16'b0000100001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000100001010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100001010101) && ({row_reg, col_reg}<16'b0000100001011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100001011001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000100001011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000100001011011) && ({row_reg, col_reg}<16'b0000100001011110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0000100001011110) && ({row_reg, col_reg}<16'b0000100001100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100001100000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000100001100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000100001100011) && ({row_reg, col_reg}<16'b0000100001101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100001101011)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b0000100001101100) && ({row_reg, col_reg}<16'b0000100001101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000100001101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000100001101111) && ({row_reg, col_reg}<16'b0000100001110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100001110001) && ({row_reg, col_reg}<16'b0000100001110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000100001110100) && ({row_reg, col_reg}<16'b0000100001110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100001110110) && ({row_reg, col_reg}<16'b0000100001111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100001111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000100001111010) && ({row_reg, col_reg}<16'b0000100010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100010000010) && ({row_reg, col_reg}<16'b0000100010101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000100010101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000100010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100010101011) && ({row_reg, col_reg}<16'b0000100010101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100010101101) && ({row_reg, col_reg}<16'b0000100010110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100010110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100010110010) && ({row_reg, col_reg}<16'b0000100010110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000100010110110) && ({row_reg, col_reg}<16'b0000100010111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000100010111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100010111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100010111010) && ({row_reg, col_reg}<16'b0000100011000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100011000100) && ({row_reg, col_reg}<16'b0000100011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000100011000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100011000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100011001000) && ({row_reg, col_reg}<16'b0000100011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100011001010) && ({row_reg, col_reg}<16'b0000100011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100011001110) && ({row_reg, col_reg}<16'b0000100011010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100011010000) && ({row_reg, col_reg}<16'b0000100011010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000100011010100) && ({row_reg, col_reg}<16'b0000100011010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100011010110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000100011010111) && ({row_reg, col_reg}<16'b0000100011011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000100011011011) && ({row_reg, col_reg}<16'b0000100011100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000100011100100) && ({row_reg, col_reg}<16'b0000100011101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100011101000) && ({row_reg, col_reg}<16'b0000100011101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000100011101011) && ({row_reg, col_reg}<16'b0000100011101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100011101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000100011101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100011101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000100011110000) && ({row_reg, col_reg}<16'b0000100011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100011110010) && ({row_reg, col_reg}<16'b0000100011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000100011111001) && ({row_reg, col_reg}<16'b0000100011111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0000100011111011) && ({row_reg, col_reg}<16'b0000100100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100100000001) && ({row_reg, col_reg}<16'b0000100100000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000100100000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100100000100) && ({row_reg, col_reg}<16'b0000100100000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100100000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100100001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100100001001) && ({row_reg, col_reg}<16'b0000100100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000100100001011) && ({row_reg, col_reg}<16'b0000100100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100100001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100100001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100100001111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0000100100010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000100100010001) && ({row_reg, col_reg}<16'b0000100100010011)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0000100100010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000100100010100) && ({row_reg, col_reg}<16'b0000100100010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000100100010111) && ({row_reg, col_reg}<16'b0000100100011001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000100100011001) && ({row_reg, col_reg}<16'b0000100100011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100100011011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000100100011100) && ({row_reg, col_reg}<16'b0000100100011111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100100011111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000100100100000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000100100100001) && ({row_reg, col_reg}<16'b0000100100100011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000100100100011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000100100100100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000100100100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000100100100110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0000100100100111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0000100100101000) && ({row_reg, col_reg}<16'b0000100100101010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000100100101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000100100101011) && ({row_reg, col_reg}<16'b0000100100101101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000100100101101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000100100101110) && ({row_reg, col_reg}<16'b0000100100110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100100110000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000100100110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000100100110010) && ({row_reg, col_reg}<16'b0000100100110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000100100110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100100110101) && ({row_reg, col_reg}<16'b0000100100110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100100110111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000100100111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100100111001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000100100111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100100111011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000100100111100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000100100111101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100100111110)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000100100111111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100101000000)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0000100101000001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0000100101000010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000100101000011) && ({row_reg, col_reg}<16'b0000100101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100101000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100101000111) && ({row_reg, col_reg}<16'b0000100101001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000100101001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000100101001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100101001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000100101001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100101001101) && ({row_reg, col_reg}<16'b0000100101001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100101001111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0000100101010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000100101010001)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}>=16'b0000100101010010) && ({row_reg, col_reg}<16'b0000100101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000100101010100) && ({row_reg, col_reg}<16'b0000100101010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100101010111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000100101011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100101011001) && ({row_reg, col_reg}<16'b0000100101011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100101011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100101011100) && ({row_reg, col_reg}<16'b0000100101011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000100101011110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000100101011111) && ({row_reg, col_reg}<16'b0000100101100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100101100001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000100101100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100101100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000100101100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100101100101) && ({row_reg, col_reg}<16'b0000100101100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000100101100111) && ({row_reg, col_reg}<16'b0000100101101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100101101001) && ({row_reg, col_reg}<16'b0000100101101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000100101101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000100101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000100101101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000100101101110) && ({row_reg, col_reg}<16'b0000100101110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000100101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100101110001) && ({row_reg, col_reg}<16'b0000100101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000100101110100) && ({row_reg, col_reg}<16'b0000100101110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100101110111) && ({row_reg, col_reg}<16'b0000100110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100110000010) && ({row_reg, col_reg}<16'b0000100110101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000100110101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000100110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100110101011) && ({row_reg, col_reg}<16'b0000100110101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100110101110) && ({row_reg, col_reg}<16'b0000100110110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100110110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100110110010) && ({row_reg, col_reg}<16'b0000100110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000100110110110) && ({row_reg, col_reg}<16'b0000100110111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000100110111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100110111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000100110111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100110111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100110111100) && ({row_reg, col_reg}<16'b0000100111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100111000101) && ({row_reg, col_reg}<16'b0000100111000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100111000111) && ({row_reg, col_reg}<16'b0000100111001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000100111001001) && ({row_reg, col_reg}<16'b0000100111001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100111001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100111001110) && ({row_reg, col_reg}<16'b0000100111010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100111010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000100111010001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000100111010010) && ({row_reg, col_reg}<16'b0000100111010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100111010101) && ({row_reg, col_reg}<16'b0000100111100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000100111100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100111100101) && ({row_reg, col_reg}<16'b0000100111100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000100111100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100111101000) && ({row_reg, col_reg}<16'b0000100111101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000100111101011) && ({row_reg, col_reg}<16'b0000100111101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100111101101) && ({row_reg, col_reg}<16'b0000100111110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000100111110000) && ({row_reg, col_reg}<16'b0000100111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100111110010) && ({row_reg, col_reg}<16'b0000100111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000100111111001) && ({row_reg, col_reg}<16'b0000100111111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0000100111111011) && ({row_reg, col_reg}<16'b0000101000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101000000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000101000000001) && ({row_reg, col_reg}<16'b0000101000000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101000000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101000000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101000000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000101000001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101000001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101000001010) && ({row_reg, col_reg}<16'b0000101000001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000101000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101000001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101000001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000101000001111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000101000010000) && ({row_reg, col_reg}<16'b0000101000010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101000010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000101000010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000101000010100) && ({row_reg, col_reg}<16'b0000101000011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000101000011000) && ({row_reg, col_reg}<16'b0000101000011010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000101000011010) && ({row_reg, col_reg}<16'b0000101000011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101000011100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000101000011101) && ({row_reg, col_reg}<16'b0000101000011111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101000011111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000101000100000) && ({row_reg, col_reg}<16'b0000101000100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101000100100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000101000100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101000100110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0000101000100111)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}>=16'b0000101000101000) && ({row_reg, col_reg}<16'b0000101000101010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000101000101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101000101011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101000101100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000101000101101) && ({row_reg, col_reg}<16'b0000101000110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101000110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000101000110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101000110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000101000110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101000110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000101000110101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0000101000110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101000110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000101000111000) && ({row_reg, col_reg}<16'b0000101000111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101000111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000101000111011) && ({row_reg, col_reg}<16'b0000101000111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101000111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101000111110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000101000111111) && ({row_reg, col_reg}<16'b0000101001000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101001000001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000101001000010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0000101001000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101001000100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0000101001000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000101001000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101001000111) && ({row_reg, col_reg}<16'b0000101001001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000101001001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000101001001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101001001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101001001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101001001111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0000101001010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000101001010001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0000101001010010)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0000101001010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000101001010100) && ({row_reg, col_reg}<16'b0000101001010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101001010110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0000101001010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000101001011000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000101001011001) && ({row_reg, col_reg}<16'b0000101001011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101001011011) && ({row_reg, col_reg}<16'b0000101001011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101001011101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0000101001011110) && ({row_reg, col_reg}<16'b0000101001100000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000101001100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000101001100001) && ({row_reg, col_reg}<16'b0000101001100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101001100011) && ({row_reg, col_reg}<16'b0000101001101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000101001101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000101001101001) && ({row_reg, col_reg}<16'b0000101001101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000101001101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000101001101100) && ({row_reg, col_reg}<16'b0000101001101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101001101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000101001101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101001110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101001110001) && ({row_reg, col_reg}<16'b0000101001110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000101001110110) && ({row_reg, col_reg}<16'b0000101001111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101001111000) && ({row_reg, col_reg}<16'b0000101001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101001111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101001111101) && ({row_reg, col_reg}<16'b0000101010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101010000011) && ({row_reg, col_reg}<16'b0000101010101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000101010101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101010101001) && ({row_reg, col_reg}<16'b0000101010101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101010101100) && ({row_reg, col_reg}<16'b0000101010101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000101010101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000101010101111) && ({row_reg, col_reg}<16'b0000101010110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101010110001) && ({row_reg, col_reg}<16'b0000101010110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000101010110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101010110111) && ({row_reg, col_reg}<16'b0000101011000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101011000110) && ({row_reg, col_reg}<16'b0000101011001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000101011001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000101011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000101011001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000101011001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000101011001101) && ({row_reg, col_reg}<16'b0000101011010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101011010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000101011010001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000101011010010) && ({row_reg, col_reg}<16'b0000101011010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000101011010100) && ({row_reg, col_reg}<16'b0000101011011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000101011011100) && ({row_reg, col_reg}<16'b0000101011100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101011100011) && ({row_reg, col_reg}<16'b0000101011100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000101011100110) && ({row_reg, col_reg}<16'b0000101011101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101011101000) && ({row_reg, col_reg}<16'b0000101011110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000101011110000) && ({row_reg, col_reg}<16'b0000101011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101011110010) && ({row_reg, col_reg}<16'b0000101011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000101011111001) && ({row_reg, col_reg}<16'b0000101011111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0000101011111011) && ({row_reg, col_reg}<16'b0000101100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101100000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000101100000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000101100000010) && ({row_reg, col_reg}<16'b0000101100000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101100000100) && ({row_reg, col_reg}<16'b0000101100000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000101100000110) && ({row_reg, col_reg}<16'b0000101100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000101100001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101100001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101100001010) && ({row_reg, col_reg}<16'b0000101100001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000101100001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000101100001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101100001110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000101100001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101100010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000101100010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101100010010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0000101100010011) && ({row_reg, col_reg}<16'b0000101100010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000101100010101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0000101100010110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000101100010111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000101100011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101100011001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000101100011010) && ({row_reg, col_reg}<16'b0000101100011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000101100011100) && ({row_reg, col_reg}<16'b0000101100011110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000101100011110) && ({row_reg, col_reg}<16'b0000101100100100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000101100100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000101100100101) && ({row_reg, col_reg}<16'b0000101100101000)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0000101100101000) && ({row_reg, col_reg}<16'b0000101100101010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000101100101010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000101100101011) && ({row_reg, col_reg}<16'b0000101100101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000101100101101) && ({row_reg, col_reg}<16'b0000101100110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101100110000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000101100110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101100110010) && ({row_reg, col_reg}<16'b0000101100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101100110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000101100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101100110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000101100111000) && ({row_reg, col_reg}<16'b0000101100111010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000101100111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000101100111011) && ({row_reg, col_reg}<16'b0000101100111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101100111101) && ({row_reg, col_reg}<16'b0000101100111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000101100111111) && ({row_reg, col_reg}<16'b0000101101000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101101000001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000101101000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101101000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000101101000100) && ({row_reg, col_reg}<16'b0000101101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000101101000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101101000111) && ({row_reg, col_reg}<16'b0000101101001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000101101001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101101001100) && ({row_reg, col_reg}<16'b0000101101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101101001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101101010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000101101010001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0000101101010010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000101101010011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000101101010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000101101010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101101010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000101101010111) && ({row_reg, col_reg}<16'b0000101101011001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000101101011001) && ({row_reg, col_reg}<16'b0000101101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101101011110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0000101101011111) && ({row_reg, col_reg}<16'b0000101101100001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000101101100001) && ({row_reg, col_reg}<16'b0000101101100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101101100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000101101100100) && ({row_reg, col_reg}<16'b0000101101101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000101101101000) && ({row_reg, col_reg}<16'b0000101101101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101101101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000101101101100) && ({row_reg, col_reg}<16'b0000101101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101101101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000101101101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101101110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101101110001) && ({row_reg, col_reg}<16'b0000101101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000101101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101101110111) && ({row_reg, col_reg}<16'b0000101101111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101101111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000101101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000101101111101) && ({row_reg, col_reg}<16'b0000101110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101110000000) && ({row_reg, col_reg}<16'b0000101110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101110000011) && ({row_reg, col_reg}<16'b0000101110101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000101110101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101110101001) && ({row_reg, col_reg}<16'b0000101110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101110101011) && ({row_reg, col_reg}<16'b0000101110101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000101110101110) && ({row_reg, col_reg}<16'b0000101110110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101110110001) && ({row_reg, col_reg}<16'b0000101110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000101110110110) && ({row_reg, col_reg}<16'b0000101111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101111000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101111000001) && ({row_reg, col_reg}<16'b0000101111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101111000111) && ({row_reg, col_reg}<16'b0000101111001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000101111001001) && ({row_reg, col_reg}<16'b0000101111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000101111001011) && ({row_reg, col_reg}<16'b0000101111001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101111001101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0000101111001110) && ({row_reg, col_reg}<16'b0000101111010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000101111010100) && ({row_reg, col_reg}<16'b0000101111010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101111010110) && ({row_reg, col_reg}<16'b0000101111011101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000101111011101) && ({row_reg, col_reg}<16'b0000101111100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101111100011) && ({row_reg, col_reg}<16'b0000101111100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000101111100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101111101000) && ({row_reg, col_reg}<16'b0000101111110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000101111110000) && ({row_reg, col_reg}<16'b0000101111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101111110010) && ({row_reg, col_reg}<16'b0000101111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000101111111001) && ({row_reg, col_reg}<16'b0000101111111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0000101111111011) && ({row_reg, col_reg}<16'b0000110000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110000000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110000000001) && ({row_reg, col_reg}<16'b0000110000000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110000000011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0000110000000100) && ({row_reg, col_reg}<16'b0000110000000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110000000110) && ({row_reg, col_reg}<16'b0000110000001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000110000001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110000001001) && ({row_reg, col_reg}<16'b0000110000001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000110000001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000110000001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000110000001111) && ({row_reg, col_reg}<16'b0000110000010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110000010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000110000010010) && ({row_reg, col_reg}<16'b0000110000010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000110000010101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0000110000010110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000110000010111) && ({row_reg, col_reg}<16'b0000110000011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000110000011001) && ({row_reg, col_reg}<16'b0000110000011011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000110000011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000110000011100) && ({row_reg, col_reg}<16'b0000110000011110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000110000011110) && ({row_reg, col_reg}<16'b0000110000100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000110000100010) && ({row_reg, col_reg}<16'b0000110000100100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000110000100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000110000100101) && ({row_reg, col_reg}<16'b0000110000101000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0000110000101000) && ({row_reg, col_reg}<16'b0000110000101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000110000101010) && ({row_reg, col_reg}<16'b0000110000101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110000101101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000110000101110) && ({row_reg, col_reg}<16'b0000110000110001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110000110001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000110000110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110000110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000110000110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000110000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110000110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000110000111000) && ({row_reg, col_reg}<16'b0000110000111010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000110000111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000110000111011) && ({row_reg, col_reg}<16'b0000110000111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000110000111101) && ({row_reg, col_reg}<16'b0000110000111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110000111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000110001000000) && ({row_reg, col_reg}<16'b0000110001000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000110001000011) && ({row_reg, col_reg}<16'b0000110001000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000110001000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110001000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110001001000) && ({row_reg, col_reg}<16'b0000110001001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000110001001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110001001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110001001101) && ({row_reg, col_reg}<16'b0000110001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110001010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000110001010001) && ({row_reg, col_reg}<16'b0000110001010011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000110001010011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000110001010100) && ({row_reg, col_reg}<16'b0000110001010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110001010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110001010111) && ({row_reg, col_reg}<16'b0000110001011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000110001011010) && ({row_reg, col_reg}<16'b0000110001011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110001011100) && ({row_reg, col_reg}<16'b0000110001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110001100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110001100011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0000110001100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000110001100101) && ({row_reg, col_reg}<16'b0000110001101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000110001101011) && ({row_reg, col_reg}<16'b0000110001101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110001101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000110001101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110001110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110001110001) && ({row_reg, col_reg}<16'b0000110001110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000110001110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110001110111) && ({row_reg, col_reg}<16'b0000110001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110001111100) && ({row_reg, col_reg}<16'b0000110001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000110001111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000110010000000) && ({row_reg, col_reg}<16'b0000110010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110010000011) && ({row_reg, col_reg}<16'b0000110010101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000110010101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000110010101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110010101010) && ({row_reg, col_reg}<16'b0000110010101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000110010101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110010101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000110010101110) && ({row_reg, col_reg}<16'b0000110010110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110010110000) && ({row_reg, col_reg}<16'b0000110010110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000110010110110) && ({row_reg, col_reg}<16'b0000110010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000110010111000) && ({row_reg, col_reg}<16'b0000110010111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110010111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000110011000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000110011000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110011000010) && ({row_reg, col_reg}<16'b0000110011000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110011000101) && ({row_reg, col_reg}<16'b0000110011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000110011001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000110011001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110011001101) && ({row_reg, col_reg}<16'b0000110011010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000110011010011) && ({row_reg, col_reg}<16'b0000110011010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110011010101) && ({row_reg, col_reg}<16'b0000110011011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000110011011100) && ({row_reg, col_reg}<16'b0000110011100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110011100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000110011100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000110011100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110011100110) && ({row_reg, col_reg}<16'b0000110011101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000110011101000) && ({row_reg, col_reg}<16'b0000110011101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110011101010) && ({row_reg, col_reg}<16'b0000110011110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000110011110000) && ({row_reg, col_reg}<16'b0000110011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110011110010) && ({row_reg, col_reg}<16'b0000110011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000110011111001) && ({row_reg, col_reg}<16'b0000110011111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0000110011111011) && ({row_reg, col_reg}<16'b0000110100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110100000000) && ({row_reg, col_reg}<16'b0000110100000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110100000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000110100000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000110100000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110100000110) && ({row_reg, col_reg}<16'b0000110100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000110100001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110100001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110100001010) && ({row_reg, col_reg}<16'b0000110100001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000110100001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110100001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110100001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110100001111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000110100010000) && ({row_reg, col_reg}<16'b0000110100010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000110100010101) && ({row_reg, col_reg}<16'b0000110100010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110100010111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000110100011000) && ({row_reg, col_reg}<16'b0000110100011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000110100011100) && ({row_reg, col_reg}<16'b0000110100011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110100011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000110100011111) && ({row_reg, col_reg}<16'b0000110100100100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110100100100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000110100100101) && ({row_reg, col_reg}<16'b0000110100101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110100101101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000110100101110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110100101111)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000110100110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110100110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110100110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000110100110011) && ({row_reg, col_reg}<16'b0000110100110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000110100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110100110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110100111000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000110100111001) && ({row_reg, col_reg}<16'b0000110100111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110100111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110100111100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000110100111101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000110100111110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000110100111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110101000000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000110101000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110101000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110101000011) && ({row_reg, col_reg}<16'b0000110101000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000110101000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110101001000) && ({row_reg, col_reg}<16'b0000110101001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000110101001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000110101001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110101001101) && ({row_reg, col_reg}<16'b0000110101001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110101001111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000110101010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110101010001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000110101010010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000110101010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110101010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110101010110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000110101010111) && ({row_reg, col_reg}<16'b0000110101011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000110101011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110101011010) && ({row_reg, col_reg}<16'b0000110101011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000110101011100) && ({row_reg, col_reg}<16'b0000110101100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110101100000) && ({row_reg, col_reg}<16'b0000110101100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110101100011) && ({row_reg, col_reg}<16'b0000110101101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000110101101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000110101101001) && ({row_reg, col_reg}<16'b0000110101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000110101101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110101101101) && ({row_reg, col_reg}<16'b0000110101101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000110101101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110101110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110101110001) && ({row_reg, col_reg}<16'b0000110101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000110101110110) && ({row_reg, col_reg}<16'b0000110101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110110000000) && ({row_reg, col_reg}<16'b0000110110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110110000011) && ({row_reg, col_reg}<16'b0000110110101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000110110101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000110110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110110101010) && ({row_reg, col_reg}<16'b0000110110101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000110110101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110110110000) && ({row_reg, col_reg}<16'b0000110110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000110110110110) && ({row_reg, col_reg}<16'b0000110110111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000110110111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000110110111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110110111011) && ({row_reg, col_reg}<16'b0000110110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110110111101) && ({row_reg, col_reg}<16'b0000110111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000110111000000) && ({row_reg, col_reg}<16'b0000110111000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110111000010) && ({row_reg, col_reg}<16'b0000110111000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110111000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000110111000101) && ({row_reg, col_reg}<16'b0000110111000111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000110111000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110111001000) && ({row_reg, col_reg}<16'b0000110111001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000110111001010) && ({row_reg, col_reg}<16'b0000110111001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000110111001110) && ({row_reg, col_reg}<16'b0000110111010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110111010000) && ({row_reg, col_reg}<16'b0000110111010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000110111010010) && ({row_reg, col_reg}<16'b0000110111010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110111010100) && ({row_reg, col_reg}<16'b0000110111011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000110111011100) && ({row_reg, col_reg}<16'b0000110111100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110111100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000110111100100) && ({row_reg, col_reg}<16'b0000110111100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110111100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000110111101000) && ({row_reg, col_reg}<16'b0000110111101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000110111101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000110111101011) && ({row_reg, col_reg}<16'b0000110111101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110111101101) && ({row_reg, col_reg}<16'b0000110111110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000110111110000) && ({row_reg, col_reg}<16'b0000110111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110111110010) && ({row_reg, col_reg}<16'b0000110111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000110111111001) && ({row_reg, col_reg}<16'b0000110111111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0000110111111011) && ({row_reg, col_reg}<16'b0000111000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111000000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000111000000001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000111000000010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111000000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000111000000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000111000000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111000000110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0000111000000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111000001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000111000001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111000001010) && ({row_reg, col_reg}<16'b0000111000001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000111000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111000001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111000001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000111000001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111000010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000111000010001)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0000111000010010) && ({row_reg, col_reg}<16'b0000111000010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000111000010110) && ({row_reg, col_reg}<16'b0000111000011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111000011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111000011001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000111000011010) && ({row_reg, col_reg}<16'b0000111000011100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000111000011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111000011101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000111000011110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000111000011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111000100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000111000100001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000111000100010) && ({row_reg, col_reg}<16'b0000111000100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000111000100101) && ({row_reg, col_reg}<16'b0000111000100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000111000100111) && ({row_reg, col_reg}<16'b0000111000101011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000111000101011) && ({row_reg, col_reg}<16'b0000111000101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111000101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111000101110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111000101111)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000111000110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111000110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111000110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000111000110011) && ({row_reg, col_reg}<16'b0000111000110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000111000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111000110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111000111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111000111001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000111000111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111000111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111000111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000111000111101) && ({row_reg, col_reg}<16'b0000111000111111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111000111111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000111001000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111001000001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000111001000010) && ({row_reg, col_reg}<16'b0000111001000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000111001000100) && ({row_reg, col_reg}<16'b0000111001000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111001000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111001001000) && ({row_reg, col_reg}<16'b0000111001001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000111001001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000111001001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111001001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111001001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111001001110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000111001001111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000111001010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111001010001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0000111001010010)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0000111001010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111001010101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000111001010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000111001010111) && ({row_reg, col_reg}<16'b0000111001011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111001011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111001011010) && ({row_reg, col_reg}<16'b0000111001011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111001011100) && ({row_reg, col_reg}<16'b0000111001100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000111001100000) && ({row_reg, col_reg}<16'b0000111001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111001100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111001100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000111001100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111001100101) && ({row_reg, col_reg}<16'b0000111001101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111001101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000111001101001) && ({row_reg, col_reg}<16'b0000111001101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000111001101011) && ({row_reg, col_reg}<16'b0000111001101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111001101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111001101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000111001101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111001110001) && ({row_reg, col_reg}<16'b0000111001110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000111001110110) && ({row_reg, col_reg}<16'b0000111001111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111001111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111001111011) && ({row_reg, col_reg}<16'b0000111010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111010000011) && ({row_reg, col_reg}<16'b0000111010101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000111010101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000111010101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111010101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000111010101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000111010101100) && ({row_reg, col_reg}<16'b0000111010101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000111010101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111010110000) && ({row_reg, col_reg}<16'b0000111010110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000111010110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000111010110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111010111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111010111001) && ({row_reg, col_reg}<16'b0000111010111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000111010111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111010111100) && ({row_reg, col_reg}<16'b0000111011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000111011000000) && ({row_reg, col_reg}<16'b0000111011000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111011000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111011000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111011000101) && ({row_reg, col_reg}<16'b0000111011001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000111011001001) && ({row_reg, col_reg}<16'b0000111011010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000111011010010) && ({row_reg, col_reg}<16'b0000111011010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111011010100) && ({row_reg, col_reg}<16'b0000111011011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111011011010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0000111011011011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000111011011100) && ({row_reg, col_reg}<16'b0000111011100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111011100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000111011100100) && ({row_reg, col_reg}<16'b0000111011100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000111011100111) && ({row_reg, col_reg}<16'b0000111011101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000111011101011) && ({row_reg, col_reg}<16'b0000111011101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000111011101101) && ({row_reg, col_reg}<16'b0000111011110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000111011110000) && ({row_reg, col_reg}<16'b0000111011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111011110010) && ({row_reg, col_reg}<16'b0000111011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000111011111001) && ({row_reg, col_reg}<16'b0000111011111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0000111011111011) && ({row_reg, col_reg}<16'b0000111100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111100000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000111100000001) && ({row_reg, col_reg}<16'b0000111100000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111100000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000111100000100) && ({row_reg, col_reg}<16'b0000111100000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111100000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000111100000111) && ({row_reg, col_reg}<16'b0000111100001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000111100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000111100001011) && ({row_reg, col_reg}<16'b0000111100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111100001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000111100001110) && ({row_reg, col_reg}<16'b0000111100010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111100010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000111100010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000111100010010) && ({row_reg, col_reg}<16'b0000111100010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000111100010110) && ({row_reg, col_reg}<16'b0000111100011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111100011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111100011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000111100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000111100011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000111100011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111100011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000111100011110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000111100011111) && ({row_reg, col_reg}<16'b0000111100100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111100100101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000111100100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111100100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000111100101000) && ({row_reg, col_reg}<16'b0000111100101010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000111100101010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000111100101011) && ({row_reg, col_reg}<16'b0000111100101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111100101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111100101110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000111100101111)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000111100110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111100110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111100110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000111100110011) && ({row_reg, col_reg}<16'b0000111100110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000111100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111100110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000111100111000) && ({row_reg, col_reg}<16'b0000111100111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111100111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111100111011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0000111100111100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000111100111101) && ({row_reg, col_reg}<16'b0000111100111111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111100111111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000111101000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111101000001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0000111101000010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000111101000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000111101000100) && ({row_reg, col_reg}<16'b0000111101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111101000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000111101000111) && ({row_reg, col_reg}<16'b0000111101001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111101001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111101001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111101001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000111101001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111101001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111101001110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0000111101001111) && ({row_reg, col_reg}<16'b0000111101010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000111101010001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0000111101010010) && ({row_reg, col_reg}<16'b0000111101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000111101010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111101010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000111101010110) && ({row_reg, col_reg}<16'b0000111101011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111101011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111101011001) && ({row_reg, col_reg}<16'b0000111101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000111101011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111101011100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000111101011101) && ({row_reg, col_reg}<16'b0000111101011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000111101011111) && ({row_reg, col_reg}<16'b0000111101100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111101100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000111101100100) && ({row_reg, col_reg}<16'b0000111101100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111101100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111101101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111101101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000111101101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000111101101011) && ({row_reg, col_reg}<16'b0000111101110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111101110001) && ({row_reg, col_reg}<16'b0000111101110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000111101110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111101110110) && ({row_reg, col_reg}<16'b0000111101111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111101111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111101111011) && ({row_reg, col_reg}<16'b0000111110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111110000011) && ({row_reg, col_reg}<16'b0000111110101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000111110101000) && ({row_reg, col_reg}<16'b0000111110101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000111110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111110101100) && ({row_reg, col_reg}<16'b0000111110101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000111110101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111110110000) && ({row_reg, col_reg}<16'b0000111110110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000111110110111) && ({row_reg, col_reg}<16'b0000111110111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111110111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000111110111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111110111100) && ({row_reg, col_reg}<16'b0000111111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111111000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000111111000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111111000010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000111111000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000111111000100) && ({row_reg, col_reg}<16'b0000111111011000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111111011000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000111111011001) && ({row_reg, col_reg}<16'b0000111111011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111111011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000111111011101) && ({row_reg, col_reg}<16'b0000111111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111111011111) && ({row_reg, col_reg}<16'b0000111111100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000111111100001) && ({row_reg, col_reg}<16'b0000111111100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111111100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000111111100100) && ({row_reg, col_reg}<16'b0000111111101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000111111101000) && ({row_reg, col_reg}<16'b0000111111101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000111111101011) && ({row_reg, col_reg}<16'b0000111111101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000111111101101) && ({row_reg, col_reg}<16'b0000111111110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000111111110000) && ({row_reg, col_reg}<16'b0000111111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111111110010) && ({row_reg, col_reg}<16'b0000111111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000111111111001) && ({row_reg, col_reg}<16'b0000111111111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0000111111111011) && ({row_reg, col_reg}<16'b0001000000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000000000000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001000000000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000000000010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001000000000011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0001000000000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000000000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000000000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000000000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000000001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001000000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001000000001010) && ({row_reg, col_reg}<16'b0001000000001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000000001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000000001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000000001111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001000000010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001000000010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000000010010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001000000010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001000000010100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0001000000010101) && ({row_reg, col_reg}<16'b0001000000010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001000000010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000000011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000000011001) && ({row_reg, col_reg}<16'b0001000000011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001000000011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001000000011100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001000000011101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001000000011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001000000011111) && ({row_reg, col_reg}<16'b0001000000100001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001000000100001) && ({row_reg, col_reg}<16'b0001000000100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000000100111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001000000101000) && ({row_reg, col_reg}<16'b0001000000101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001000000101010) && ({row_reg, col_reg}<16'b0001000000101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000000101100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001000000101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000000101110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001000000101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001000000110000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001000000110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000000110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001000000110011) && ({row_reg, col_reg}<16'b0001000000110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001000000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000000110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000000111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001000000111001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001000000111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000000111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000000111100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001000000111101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001000000111110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001000000111111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001000001000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000001000001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0001000001000010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001000001000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000001000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000001000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000001000110) && ({row_reg, col_reg}<16'b0001000001001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000001001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001000001001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001000001001101) && ({row_reg, col_reg}<16'b0001000001001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001000001001111) && ({row_reg, col_reg}<16'b0001000001010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001000001010011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0001000001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000001010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000001010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000001010111) && ({row_reg, col_reg}<16'b0001000001011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001000001011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000001011100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001000001011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001000001011110) && ({row_reg, col_reg}<16'b0001000001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000001100010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001000001100011) && ({row_reg, col_reg}<16'b0001000001100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000001100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001000001101000) && ({row_reg, col_reg}<16'b0001000001101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001000001101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001000001101011) && ({row_reg, col_reg}<16'b0001000001101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000001101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001000001101111) && ({row_reg, col_reg}<16'b0001000001110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000001110001) && ({row_reg, col_reg}<16'b0001000001110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001000001110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000001110110) && ({row_reg, col_reg}<16'b0001000010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000010000011) && ({row_reg, col_reg}<16'b0001000010101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001000010101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001000010101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001000010101011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=16'b0001000010101100) && ({row_reg, col_reg}<16'b0001000010101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001000010101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000010110000) && ({row_reg, col_reg}<16'b0001000010110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001000010110110) && ({row_reg, col_reg}<16'b0001000010111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000010111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000010111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001000010111110) && ({row_reg, col_reg}<16'b0001000011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000011000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001000011000001) && ({row_reg, col_reg}<16'b0001000011000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000011000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000011000100) && ({row_reg, col_reg}<16'b0001000011001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001000011001011) && ({row_reg, col_reg}<16'b0001000011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000011001110) && ({row_reg, col_reg}<16'b0001000011010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000011010010) && ({row_reg, col_reg}<16'b0001000011010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000011010101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001000011010110) && ({row_reg, col_reg}<16'b0001000011011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000011011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001000011011101) && ({row_reg, col_reg}<16'b0001000011100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000011100000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001000011100001) && ({row_reg, col_reg}<16'b0001000011100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000011100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001000011100100) && ({row_reg, col_reg}<16'b0001000011101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001000011101000) && ({row_reg, col_reg}<16'b0001000011101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001000011101011) && ({row_reg, col_reg}<16'b0001000011101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001000011101101) && ({row_reg, col_reg}<16'b0001000011110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001000011110000) && ({row_reg, col_reg}<16'b0001000011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000011110010) && ({row_reg, col_reg}<16'b0001000011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001000011111001) && ({row_reg, col_reg}<16'b0001000011111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0001000011111011) && ({row_reg, col_reg}<16'b0001000100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000100000000) && ({row_reg, col_reg}<16'b0001000100000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001000100000010) && ({row_reg, col_reg}<16'b0001000100000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000100000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000100000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001000100001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000100001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001000100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000100001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000100001100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001000100001101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0001000100001110) && ({row_reg, col_reg}<16'b0001000100010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001000100010000) && ({row_reg, col_reg}<16'b0001000100010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000100010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001000100010011) && ({row_reg, col_reg}<16'b0001000100010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001000100010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000100010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001000100010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000100011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000100011001) && ({row_reg, col_reg}<16'b0001000100011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001000100011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000100011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000100011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001000100011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001000100011111) && ({row_reg, col_reg}<16'b0001000100100001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001000100100001) && ({row_reg, col_reg}<16'b0001000100100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001000100100110) && ({row_reg, col_reg}<16'b0001000100101000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001000100101000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0001000100101001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001000100101010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001000100101011) && ({row_reg, col_reg}<16'b0001000100101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000100101110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001000100101111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001000100110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001000100110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000100110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001000100110011) && ({row_reg, col_reg}<16'b0001000100110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001000100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000100110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000100111000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001000100111001) && ({row_reg, col_reg}<16'b0001000100111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001000100111011) && ({row_reg, col_reg}<16'b0001000100111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001000100111101) && ({row_reg, col_reg}<16'b0001000101000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001000101000001) && ({row_reg, col_reg}<16'b0001000101000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001000101000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000101000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000101000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000101000110) && ({row_reg, col_reg}<16'b0001000101001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000101001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001000101001011) && ({row_reg, col_reg}<16'b0001000101001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000101001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001000101001110) && ({row_reg, col_reg}<16'b0001000101010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000101010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001000101010001) && ({row_reg, col_reg}<16'b0001000101010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001000101010011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0001000101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000101010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000101010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000101010111) && ({row_reg, col_reg}<16'b0001000101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001000101011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000101011100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001000101011101) && ({row_reg, col_reg}<16'b0001000101100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000101100010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001000101100011) && ({row_reg, col_reg}<16'b0001000101100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000101100110) && ({row_reg, col_reg}<16'b0001000101101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001000101101001) && ({row_reg, col_reg}<16'b0001000101101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000101101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001000101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000101101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001000101101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000101101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000101110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000101110001) && ({row_reg, col_reg}<16'b0001000101110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001000101110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000101110110) && ({row_reg, col_reg}<16'b0001000101111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000101111001) && ({row_reg, col_reg}<16'b0001000101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000101111011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==16'b0001000101111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000101111101) && ({row_reg, col_reg}<16'b0001000101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000101111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001000110000000) && ({row_reg, col_reg}<16'b0001000110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000110000011) && ({row_reg, col_reg}<16'b0001000110101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001000110101000) && ({row_reg, col_reg}<16'b0001000110101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001000110101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000110110000) && ({row_reg, col_reg}<16'b0001000110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001000110110110) && ({row_reg, col_reg}<16'b0001000110111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000110111011) && ({row_reg, col_reg}<16'b0001000110111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001000110111101) && ({row_reg, col_reg}<16'b0001000110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001000110111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000111000001) && ({row_reg, col_reg}<16'b0001000111000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000111000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000111000101) && ({row_reg, col_reg}<16'b0001000111001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000111001001) && ({row_reg, col_reg}<16'b0001000111001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001000111001011) && ({row_reg, col_reg}<16'b0001000111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000111001110) && ({row_reg, col_reg}<16'b0001000111010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000111010010) && ({row_reg, col_reg}<16'b0001000111010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001000111010101) && ({row_reg, col_reg}<16'b0001000111010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000111010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001000111011000) && ({row_reg, col_reg}<16'b0001000111011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000111011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001000111011101) && ({row_reg, col_reg}<16'b0001000111100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000111100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000111100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000111100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001000111100100) && ({row_reg, col_reg}<16'b0001000111101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001000111101000) && ({row_reg, col_reg}<16'b0001000111101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001000111101011) && ({row_reg, col_reg}<16'b0001000111101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001000111101101) && ({row_reg, col_reg}<16'b0001000111110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001000111110000) && ({row_reg, col_reg}<16'b0001000111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000111110010) && ({row_reg, col_reg}<16'b0001000111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001000111111001) && ({row_reg, col_reg}<16'b0001000111111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0001000111111011) && ({row_reg, col_reg}<16'b0001001000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001000000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001000000001) && ({row_reg, col_reg}<16'b0001001000000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001001000000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001000000100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0001001000000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001000000110) && ({row_reg, col_reg}<16'b0001001000001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001000001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001001000001001) && ({row_reg, col_reg}<16'b0001001000001100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001001000001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001000001101) && ({row_reg, col_reg}<16'b0001001000010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001001000010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001000010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001000010010) && ({row_reg, col_reg}<16'b0001001000010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001001000010100) && ({row_reg, col_reg}<16'b0001001000010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001001000010110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0001001000010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001000011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001000011001) && ({row_reg, col_reg}<16'b0001001000011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001001000011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001000011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001000011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001001000011110) && ({row_reg, col_reg}<16'b0001001000100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001001000100110) && ({row_reg, col_reg}<16'b0001001000101000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001001000101000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0001001000101001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001001000101010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001001000101011) && ({row_reg, col_reg}<16'b0001001000101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001001000101110) && ({row_reg, col_reg}<16'b0001001000110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001001000110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001001000110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001001000110010) && ({row_reg, col_reg}<16'b0001001000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001000110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001000110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001000110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001001000111000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001001000111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001001000111010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001001000111011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0001001000111100) && ({row_reg, col_reg}<16'b0001001001000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001001001000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001001001000100) && ({row_reg, col_reg}<16'b0001001001000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001001000110) && ({row_reg, col_reg}<16'b0001001001001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001001001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001001001001011) && ({row_reg, col_reg}<16'b0001001001001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001001001001101) && ({row_reg, col_reg}<16'b0001001001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001001001111) && ({row_reg, col_reg}<16'b0001001001010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001001001010001) && ({row_reg, col_reg}<16'b0001001001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001001001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001001010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001001010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001001010111) && ({row_reg, col_reg}<16'b0001001001011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001001001011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001001011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001001011101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0001001001011110) && ({row_reg, col_reg}<16'b0001001001100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001001100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001001100010) && ({row_reg, col_reg}<16'b0001001001100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001001001100100) && ({row_reg, col_reg}<16'b0001001001100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001001001100110) && ({row_reg, col_reg}<16'b0001001001101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001001001101001) && ({row_reg, col_reg}<16'b0001001001101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001001101011) && ({row_reg, col_reg}<16'b0001001001101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001001001101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001001110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001001110001) && ({row_reg, col_reg}<16'b0001001001110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001001001110110) && ({row_reg, col_reg}<16'b0001001001111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001001111001) && ({row_reg, col_reg}<16'b0001001001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001001111011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==16'b0001001001111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001001001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001001001111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001001010000000) && ({row_reg, col_reg}<16'b0001001010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001010000011) && ({row_reg, col_reg}<16'b0001001010101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001001010101000) && ({row_reg, col_reg}<16'b0001001010101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001010101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001001010101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001001010101101) && ({row_reg, col_reg}<16'b0001001010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001001010110000) && ({row_reg, col_reg}<16'b0001001010110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001001010110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001010110110) && ({row_reg, col_reg}<16'b0001001010111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001010111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001001010111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001010111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001001010111101) && ({row_reg, col_reg}<16'b0001001011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001011000001) && ({row_reg, col_reg}<16'b0001001011000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001011000100) && ({row_reg, col_reg}<16'b0001001011000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001011000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001001011001000) && ({row_reg, col_reg}<16'b0001001011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001011001010) && ({row_reg, col_reg}<16'b0001001011001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001011001100) && ({row_reg, col_reg}<16'b0001001011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001011001110) && ({row_reg, col_reg}<16'b0001001011010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001011010101) && ({row_reg, col_reg}<16'b0001001011011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001011011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001011011101) && ({row_reg, col_reg}<16'b0001001011100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001011100001) && ({row_reg, col_reg}<16'b0001001011100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001011100100) && ({row_reg, col_reg}<16'b0001001011100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001011100111) && ({row_reg, col_reg}<16'b0001001011101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001001011101010) && ({row_reg, col_reg}<16'b0001001011101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001011101101) && ({row_reg, col_reg}<16'b0001001011110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001011110000) && ({row_reg, col_reg}<16'b0001001011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001011110010) && ({row_reg, col_reg}<16'b0001001011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001001011111001) && ({row_reg, col_reg}<16'b0001001011111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0001001011111011) && ({row_reg, col_reg}<16'b0001001100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001100000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001001100000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001100000010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001001100000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001100000100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0001001100000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001100000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001001100000111) && ({row_reg, col_reg}<16'b0001001100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001001100001010) && ({row_reg, col_reg}<16'b0001001100001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001100001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001100001101) && ({row_reg, col_reg}<16'b0001001100010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001001100010000) && ({row_reg, col_reg}<16'b0001001100010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001100010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001001100010011) && ({row_reg, col_reg}<16'b0001001100010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001001100010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001100010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001100011000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001100011001) && ({row_reg, col_reg}<16'b0001001100011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001100011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001100011101) && ({row_reg, col_reg}<16'b0001001100011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001100011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001001100100000) && ({row_reg, col_reg}<16'b0001001100100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001001100100101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001001100100110) && ({row_reg, col_reg}<16'b0001001100101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001001100101010)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0001001100101011) && ({row_reg, col_reg}<16'b0001001100101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001001100101110) && ({row_reg, col_reg}<16'b0001001100110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001001100110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001001100110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001001100110010) && ({row_reg, col_reg}<16'b0001001100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001100110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001100110101) && ({row_reg, col_reg}<16'b0001001100110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001100110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001001100111000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001001100111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001001100111010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001001100111011)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0001001100111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001001100111101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001001100111110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0001001100111111) && ({row_reg, col_reg}<16'b0001001101000001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001001101000001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0001001101000010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001001101000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001001101000100) && ({row_reg, col_reg}<16'b0001001101001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001101001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001101001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001101001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001001101001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001001101001100) && ({row_reg, col_reg}<16'b0001001101010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001101010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001001101010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001001101010010)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0001001101010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001001101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001101010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001101010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001101010111) && ({row_reg, col_reg}<16'b0001001101011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001101011001) && ({row_reg, col_reg}<16'b0001001101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001001101011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001101011100) && ({row_reg, col_reg}<16'b0001001101011110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001101011110) && ({row_reg, col_reg}<16'b0001001101100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001101100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001001101100100) && ({row_reg, col_reg}<16'b0001001101100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001001101100111) && ({row_reg, col_reg}<16'b0001001101101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001001101101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001101101010) && ({row_reg, col_reg}<16'b0001001101101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001001101101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001101110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001101110001) && ({row_reg, col_reg}<16'b0001001101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001001101110110) && ({row_reg, col_reg}<16'b0001001101111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001101111001) && ({row_reg, col_reg}<16'b0001001101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001101111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001001101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001001101111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001001101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001001101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001110000000) && ({row_reg, col_reg}<16'b0001001110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001110000011) && ({row_reg, col_reg}<16'b0001001110101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001001110101000) && ({row_reg, col_reg}<16'b0001001110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001110101101) && ({row_reg, col_reg}<16'b0001001110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001110110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001110110001) && ({row_reg, col_reg}<16'b0001001110110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001001110110101) && ({row_reg, col_reg}<16'b0001001110111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001110111000) && ({row_reg, col_reg}<16'b0001001110111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001001110111010) && ({row_reg, col_reg}<16'b0001001110111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001110111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001001110111101) && ({row_reg, col_reg}<16'b0001001111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001001111000000) && ({row_reg, col_reg}<16'b0001001111000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001111000011) && ({row_reg, col_reg}<16'b0001001111000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001111000110) && ({row_reg, col_reg}<16'b0001001111001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001001111001010) && ({row_reg, col_reg}<16'b0001001111010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001111010010) && ({row_reg, col_reg}<16'b0001001111010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001111010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001111010101) && ({row_reg, col_reg}<16'b0001001111011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001111011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001111011101) && ({row_reg, col_reg}<16'b0001001111100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001111100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001111100100) && ({row_reg, col_reg}<16'b0001001111101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001111101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001111101110) && ({row_reg, col_reg}<16'b0001001111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001111110010) && ({row_reg, col_reg}<16'b0001001111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001001111111001) && ({row_reg, col_reg}<16'b0001001111111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0001001111111011) && ({row_reg, col_reg}<16'b0001010000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010000000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001010000000001) && ({row_reg, col_reg}<16'b0001010000000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010000000100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0001010000000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001010000000110) && ({row_reg, col_reg}<16'b0001010000001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010000001100) && ({row_reg, col_reg}<16'b0001010000001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010000001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010000001111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001010000010000) && ({row_reg, col_reg}<16'b0001010000010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010000010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010000010011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001010000010100) && ({row_reg, col_reg}<16'b0001010000010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010000010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001010000010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010000011000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001010000011001) && ({row_reg, col_reg}<16'b0001010000011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010000011011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010000011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010000011101) && ({row_reg, col_reg}<16'b0001010000011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010000011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001010000100000) && ({row_reg, col_reg}<16'b0001010000100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010000100100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001010000100101) && ({row_reg, col_reg}<16'b0001010000101000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010000101000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0001010000101001) && ({row_reg, col_reg}<16'b0001010000101011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0001010000101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001010000101100) && ({row_reg, col_reg}<16'b0001010000101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001010000101110) && ({row_reg, col_reg}<16'b0001010000110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001010000110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010000110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001010000110010) && ({row_reg, col_reg}<16'b0001010000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010000110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010000110101) && ({row_reg, col_reg}<16'b0001010000110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010000110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010000111000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001010000111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010000111010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001010000111011) && ({row_reg, col_reg}<16'b0001010000111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010000111101) && ({row_reg, col_reg}<16'b0001010001000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010001000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001010001000001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0001010001000010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001010001000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010001000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010001000101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001010001000110) && ({row_reg, col_reg}<16'b0001010001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010001001001) && ({row_reg, col_reg}<16'b0001010001001100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001010001001100) && ({row_reg, col_reg}<16'b0001010001010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010001010000) && ({row_reg, col_reg}<16'b0001010001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001010001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010001010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001010001010110) && ({row_reg, col_reg}<16'b0001010001011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010001011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001010001011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001010001011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010001011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010001011101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0001010001011110) && ({row_reg, col_reg}<16'b0001010001100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010001100100) && ({row_reg, col_reg}<16'b0001010001101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010001101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001010001101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010001101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010001101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001010001101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010001101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010001101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001010001101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010001110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010001110001) && ({row_reg, col_reg}<16'b0001010001110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001010001110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010001110111) && ({row_reg, col_reg}<16'b0001010001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010001111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001010001111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001010001111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001010001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010010000000) && ({row_reg, col_reg}<16'b0001010010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010010000011) && ({row_reg, col_reg}<16'b0001010010101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001010010101000) && ({row_reg, col_reg}<16'b0001010010101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010010101100) && ({row_reg, col_reg}<16'b0001010010101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001010010101111) && ({row_reg, col_reg}<16'b0001010010110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010010110001) && ({row_reg, col_reg}<16'b0001010010110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001010010110101) && ({row_reg, col_reg}<16'b0001010010111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010010111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010010111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010010111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001010010111011) && ({row_reg, col_reg}<16'b0001010010111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010010111101) && ({row_reg, col_reg}<16'b0001010011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001010011000000) && ({row_reg, col_reg}<16'b0001010011000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010011000101) && ({row_reg, col_reg}<16'b0001010011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001010011001011) && ({row_reg, col_reg}<16'b0001010011010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001010011010010) && ({row_reg, col_reg}<16'b0001010011010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010011010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010011010101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001010011010110) && ({row_reg, col_reg}<16'b0001010011011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010011011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001010011011101) && ({row_reg, col_reg}<16'b0001010011100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010011100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001010011100100) && ({row_reg, col_reg}<16'b0001010011101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010011101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001010011101110) && ({row_reg, col_reg}<16'b0001010011110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010011110010) && ({row_reg, col_reg}<16'b0001010011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001010011111001) && ({row_reg, col_reg}<16'b0001010011111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0001010011111011) && ({row_reg, col_reg}<16'b0001010100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010100000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001010100000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001010100000010) && ({row_reg, col_reg}<16'b0001010100000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010100000101) && ({row_reg, col_reg}<16'b0001010100000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001010100001000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001010100001001)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0001010100001010) && ({row_reg, col_reg}<16'b0001010100001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010100001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010100001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001010100001110) && ({row_reg, col_reg}<16'b0001010100010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001010100010000) && ({row_reg, col_reg}<16'b0001010100010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010100010010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001010100010011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001010100010100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001010100010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010100010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001010100010111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0001010100011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010100011001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001010100011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010100011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001010100011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010100011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010100011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001010100011111) && ({row_reg, col_reg}<16'b0001010100100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010100100100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001010100100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010100100110)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0001010100100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001010100101000) && ({row_reg, col_reg}<16'b0001010100101010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0001010100101010)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0001010100101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001010100101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001010100101101) && ({row_reg, col_reg}<16'b0001010100101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001010100101111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001010100110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010100110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001010100110010) && ({row_reg, col_reg}<16'b0001010100110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010100110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010100110101) && ({row_reg, col_reg}<16'b0001010100110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010100110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010100111000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001010100111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010100111010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001010100111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010100111100) && ({row_reg, col_reg}<16'b0001010100111110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001010100111110) && ({row_reg, col_reg}<16'b0001010101000000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001010101000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010101000001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001010101000010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0001010101000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010101000100)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}>=16'b0001010101000101) && ({row_reg, col_reg}<16'b0001010101000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010101000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001010101001000) && ({row_reg, col_reg}<16'b0001010101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010101001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001010101001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010101001101) && ({row_reg, col_reg}<16'b0001010101001111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0001010101001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010101010000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0001010101010001) && ({row_reg, col_reg}<16'b0001010101010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010101010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010101010110) && ({row_reg, col_reg}<16'b0001010101011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001010101011001) && ({row_reg, col_reg}<16'b0001010101011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001010101011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010101011100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0001010101011101) && ({row_reg, col_reg}<16'b0001010101011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001010101011111) && ({row_reg, col_reg}<16'b0001010101100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010101100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001010101100100)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b0001010101100101) && ({row_reg, col_reg}<16'b0001010101101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010101101001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001010101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010101101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010101101100) && ({row_reg, col_reg}<16'b0001010101101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010101101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010101110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010101110001) && ({row_reg, col_reg}<16'b0001010101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001010101110110) && ({row_reg, col_reg}<16'b0001010101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010101111000) && ({row_reg, col_reg}<16'b0001010101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010101111100) && ({row_reg, col_reg}<16'b0001010110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010110000000) && ({row_reg, col_reg}<16'b0001010110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010110000011) && ({row_reg, col_reg}<16'b0001010110101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001010110101000) && ({row_reg, col_reg}<16'b0001010110101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010110101100) && ({row_reg, col_reg}<16'b0001010110101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001010110101111) && ({row_reg, col_reg}<16'b0001010110110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010110110001) && ({row_reg, col_reg}<16'b0001010110110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001010110110101) && ({row_reg, col_reg}<16'b0001010110110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010110110111) && ({row_reg, col_reg}<16'b0001010110111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010110111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010110111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001010110111011) && ({row_reg, col_reg}<16'b0001010110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010110111101) && ({row_reg, col_reg}<16'b0001010111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001010111000000) && ({row_reg, col_reg}<16'b0001010111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010111000101) && ({row_reg, col_reg}<16'b0001010111001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010111001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010111001101) && ({row_reg, col_reg}<16'b0001010111010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010111010101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001010111010110) && ({row_reg, col_reg}<16'b0001010111011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010111011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001010111011101) && ({row_reg, col_reg}<16'b0001010111100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010111100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010111100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010111100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001010111100100) && ({row_reg, col_reg}<16'b0001010111101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010111101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001010111101001) && ({row_reg, col_reg}<16'b0001010111101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010111101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001010111101110) && ({row_reg, col_reg}<16'b0001010111110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010111110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010111110010) && ({row_reg, col_reg}<16'b0001010111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001010111111001) && ({row_reg, col_reg}<16'b0001010111111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0001010111111011) && ({row_reg, col_reg}<16'b0001011000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011000000000) && ({row_reg, col_reg}<16'b0001011000000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011000000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011000000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001011000000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011000000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011000000110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0001011000000111) && ({row_reg, col_reg}<16'b0001011000001010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001011000001010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0001011000001011) && ({row_reg, col_reg}<16'b0001011000001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011000001101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001011000001110) && ({row_reg, col_reg}<16'b0001011000010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011000010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011000010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001011000010010) && ({row_reg, col_reg}<16'b0001011000010100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001011000010100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001011000010101) && ({row_reg, col_reg}<16'b0001011000011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011000011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011000011001) && ({row_reg, col_reg}<16'b0001011000011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011000011100) && ({row_reg, col_reg}<16'b0001011000011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011000011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001011000011111) && ({row_reg, col_reg}<16'b0001011000100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011000100101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001011000100110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001011000100111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001011000101000)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0001011000101001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0001011000101010) && ({row_reg, col_reg}<16'b0001011000101100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001011000101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011000101101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001011000101110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001011000101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001011000110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011000110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011000110010) && ({row_reg, col_reg}<16'b0001011000110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001011000110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011000110101) && ({row_reg, col_reg}<16'b0001011000110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011000110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011000111000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001011000111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011000111010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001011000111011) && ({row_reg, col_reg}<16'b0001011000111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011000111101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001011000111110) && ({row_reg, col_reg}<16'b0001011001000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011001000001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001011001000010) && ({row_reg, col_reg}<16'b0001011001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011001000110) && ({row_reg, col_reg}<16'b0001011001001000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001011001001000) && ({row_reg, col_reg}<16'b0001011001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011001001010) && ({row_reg, col_reg}<16'b0001011001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011001001110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0001011001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011001010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001011001010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001011001010010) && ({row_reg, col_reg}<16'b0001011001010100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001011001010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001011001010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011001010110) && ({row_reg, col_reg}<16'b0001011001011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001011001011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011001011010) && ({row_reg, col_reg}<16'b0001011001011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011001011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011001011101) && ({row_reg, col_reg}<16'b0001011001100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011001100000) && ({row_reg, col_reg}<16'b0001011001100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011001100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001011001100100)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b0001011001100101) && ({row_reg, col_reg}<16'b0001011001101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011001101011) && ({row_reg, col_reg}<16'b0001011001101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011001101101) && ({row_reg, col_reg}<16'b0001011001110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001011001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011001110001) && ({row_reg, col_reg}<16'b0001011001110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001011001110110) && ({row_reg, col_reg}<16'b0001011001111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011001111001) && ({row_reg, col_reg}<16'b0001011001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001011001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011001111100) && ({row_reg, col_reg}<16'b0001011010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011010000000) && ({row_reg, col_reg}<16'b0001011010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011010000011) && ({row_reg, col_reg}<16'b0001011010100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001011010100111) && ({row_reg, col_reg}<16'b0001011010101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011010101001) && ({row_reg, col_reg}<16'b0001011010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011010101101) && ({row_reg, col_reg}<16'b0001011010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001011010110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011010110001) && ({row_reg, col_reg}<16'b0001011010110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001011010110101) && ({row_reg, col_reg}<16'b0001011010111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011010111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001011010111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011010111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001011010111011) && ({row_reg, col_reg}<16'b0001011010111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011010111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001011010111110) && ({row_reg, col_reg}<16'b0001011011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011011000000) && ({row_reg, col_reg}<16'b0001011011000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011011000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011011000110) && ({row_reg, col_reg}<16'b0001011011001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001011011001000) && ({row_reg, col_reg}<16'b0001011011001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001011011001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011011001110) && ({row_reg, col_reg}<16'b0001011011010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001011011010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011011010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001011011010101) && ({row_reg, col_reg}<16'b0001011011011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011011011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011011011010) && ({row_reg, col_reg}<16'b0001011011011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011011011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001011011011101) && ({row_reg, col_reg}<16'b0001011011100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011011100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001011011100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011011100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001011011100100) && ({row_reg, col_reg}<16'b0001011011101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011011101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011011101011) && ({row_reg, col_reg}<16'b0001011011101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011011101101) && ({row_reg, col_reg}<16'b0001011011101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001011011101111) && ({row_reg, col_reg}<16'b0001011011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011011110010) && ({row_reg, col_reg}<16'b0001011011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001011011111001) && ({row_reg, col_reg}<16'b0001011011111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0001011011111011) && ({row_reg, col_reg}<16'b0001011100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011100000000) && ({row_reg, col_reg}<16'b0001011100000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011100000010) && ({row_reg, col_reg}<16'b0001011100000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001011100000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011100000110) && ({row_reg, col_reg}<16'b0001011100001000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001011100001000) && ({row_reg, col_reg}<16'b0001011100001010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0001011100001010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011100001011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001011100001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011100001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001011100001110) && ({row_reg, col_reg}<16'b0001011100010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011100010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001011100010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011100010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001011100010011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0001011100010100) && ({row_reg, col_reg}<16'b0001011100010110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001011100010110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001011100010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011100011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011100011001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0001011100011010) && ({row_reg, col_reg}<16'b0001011100011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001011100011100) && ({row_reg, col_reg}<16'b0001011100011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011100011110) && ({row_reg, col_reg}<16'b0001011100101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011100101001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001011100101010) && ({row_reg, col_reg}<16'b0001011100101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011100101100) && ({row_reg, col_reg}<16'b0001011100101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001011100101110) && ({row_reg, col_reg}<16'b0001011100110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001011100110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011100110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011100110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011100110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011100110100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001011100110101)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0001011100110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011100110111) && ({row_reg, col_reg}<16'b0001011100111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011100111010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001011100111011) && ({row_reg, col_reg}<16'b0001011100111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011100111101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001011100111110) && ({row_reg, col_reg}<16'b0001011101000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011101000001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001011101000010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0001011101000011) && ({row_reg, col_reg}<16'b0001011101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011101000110) && ({row_reg, col_reg}<16'b0001011101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001011101001001) && ({row_reg, col_reg}<16'b0001011101001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011101001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011101001110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0001011101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011101010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001011101010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011101010010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001011101010011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001011101010100) && ({row_reg, col_reg}<16'b0001011101010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011101010110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001011101010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011101011000) && ({row_reg, col_reg}<16'b0001011101011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011101011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001011101011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011101011101) && ({row_reg, col_reg}<16'b0001011101100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011101100000) && ({row_reg, col_reg}<16'b0001011101100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011101100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001011101100100) && ({row_reg, col_reg}<16'b0001011101100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001011101100110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001011101100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001011101101000) && ({row_reg, col_reg}<16'b0001011101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011101101010) && ({row_reg, col_reg}<16'b0001011101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011101101110) && ({row_reg, col_reg}<16'b0001011101110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001011101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011101110001) && ({row_reg, col_reg}<16'b0001011101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001011101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011101110111) && ({row_reg, col_reg}<16'b0001011101111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011101111001) && ({row_reg, col_reg}<16'b0001011101111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011101111100) && ({row_reg, col_reg}<16'b0001011110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011110000000) && ({row_reg, col_reg}<16'b0001011110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011110000011) && ({row_reg, col_reg}<16'b0001011110100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001011110100100) && ({row_reg, col_reg}<16'b0001011110100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011110100110) && ({row_reg, col_reg}<16'b0001011110101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011110101000) && ({row_reg, col_reg}<16'b0001011110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011110101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011110101011) && ({row_reg, col_reg}<16'b0001011110101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001011110101110) && ({row_reg, col_reg}<16'b0001011110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011110110000) && ({row_reg, col_reg}<16'b0001011110110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001011110110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011110110101) && ({row_reg, col_reg}<16'b0001011110110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011110110111) && ({row_reg, col_reg}<16'b0001011110111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001011110111011) && ({row_reg, col_reg}<16'b0001011110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011110111101) && ({row_reg, col_reg}<16'b0001011110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001011110111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011111000000) && ({row_reg, col_reg}<16'b0001011111000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011111000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011111000101) && ({row_reg, col_reg}<16'b0001011111001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001011111001001) && ({row_reg, col_reg}<16'b0001011111001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011111001101) && ({row_reg, col_reg}<16'b0001011111010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001011111010010) && ({row_reg, col_reg}<16'b0001011111010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011111010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001011111010101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0001011111010110) && ({row_reg, col_reg}<16'b0001011111011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011111011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001011111011101) && ({row_reg, col_reg}<16'b0001011111100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011111100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001011111100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011111100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001011111100100) && ({row_reg, col_reg}<16'b0001011111101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011111101101) && ({row_reg, col_reg}<16'b0001011111110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001011111110000) && ({row_reg, col_reg}<16'b0001011111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011111110010) && ({row_reg, col_reg}<16'b0001011111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001011111111001) && ({row_reg, col_reg}<16'b0001011111111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0001011111111011) && ({row_reg, col_reg}<16'b0001100000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100000000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100000000001) && ({row_reg, col_reg}<16'b0001100000000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001100000000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001100000000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100000000110) && ({row_reg, col_reg}<16'b0001100000001000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001100000001000) && ({row_reg, col_reg}<16'b0001100000001010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001100000001010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100000001011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001100000001100) && ({row_reg, col_reg}<16'b0001100000010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100000010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100000010010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0001100000010011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0001100000010100)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0001100000010101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0001100000010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100000010111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001100000011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100000011001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001100000011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001100000011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100000011100) && ({row_reg, col_reg}<16'b0001100000011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100000011110) && ({row_reg, col_reg}<16'b0001100000100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001100000100001) && ({row_reg, col_reg}<16'b0001100000100011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001100000100011) && ({row_reg, col_reg}<16'b0001100000100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100000100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001100000100110)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0001100000100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001100000101000) && ({row_reg, col_reg}<16'b0001100000101010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001100000101010) && ({row_reg, col_reg}<16'b0001100000101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100000101100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001100000101101) && ({row_reg, col_reg}<16'b0001100000110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001100000110001) && ({row_reg, col_reg}<16'b0001100000110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100000110011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0001100000110100) && ({row_reg, col_reg}<16'b0001100000111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100000111001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001100000111010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0001100000111011) && ({row_reg, col_reg}<16'b0001100000111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100000111101) && ({row_reg, col_reg}<16'b0001100000111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100000111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001100001000000) && ({row_reg, col_reg}<16'b0001100001000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001100001000011) && ({row_reg, col_reg}<16'b0001100001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100001000110) && ({row_reg, col_reg}<16'b0001100001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100001001001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001100001001010) && ({row_reg, col_reg}<16'b0001100001001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100001001110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0001100001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100001010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001100001010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100001010010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001100001010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001100001010100) && ({row_reg, col_reg}<16'b0001100001010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100001010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100001010111) && ({row_reg, col_reg}<16'b0001100001011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100001011010) && ({row_reg, col_reg}<16'b0001100001011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001100001011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100001011101) && ({row_reg, col_reg}<16'b0001100001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100001011111) && ({row_reg, col_reg}<16'b0001100001100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100001100010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0001100001100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001100001100100) && ({row_reg, col_reg}<16'b0001100001100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100001100110) && ({row_reg, col_reg}<16'b0001100001101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001100001101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100001101001) && ({row_reg, col_reg}<16'b0001100001101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100001101101) && ({row_reg, col_reg}<16'b0001100001110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001100001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100001110001) && ({row_reg, col_reg}<16'b0001100001110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100001110011) && ({row_reg, col_reg}<16'b0001100001110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001100001110101) && ({row_reg, col_reg}<16'b0001100001111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001100001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100001111001) && ({row_reg, col_reg}<16'b0001100001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001100001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100001111100) && ({row_reg, col_reg}<16'b0001100001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100001111110) && ({row_reg, col_reg}<16'b0001100010000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001100010000000) && ({row_reg, col_reg}<16'b0001100010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100010000011) && ({row_reg, col_reg}<16'b0001100010100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001100010100011) && ({row_reg, col_reg}<16'b0001100010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100010101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100010101011) && ({row_reg, col_reg}<16'b0001100010101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001100010101110) && ({row_reg, col_reg}<16'b0001100010110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100010110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100010110001) && ({row_reg, col_reg}<16'b0001100010110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001100010110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100010110101) && ({row_reg, col_reg}<16'b0001100010110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100010110111) && ({row_reg, col_reg}<16'b0001100010111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001100010111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001100010111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100010111101) && ({row_reg, col_reg}<16'b0001100010111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001100010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100011000000) && ({row_reg, col_reg}<16'b0001100011000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100011000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100011000101) && ({row_reg, col_reg}<16'b0001100011001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001100011001001) && ({row_reg, col_reg}<16'b0001100011001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100011001101) && ({row_reg, col_reg}<16'b0001100011010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001100011010010) && ({row_reg, col_reg}<16'b0001100011010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100011010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001100011010101) && ({row_reg, col_reg}<16'b0001100011011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100011011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001100011011101) && ({row_reg, col_reg}<16'b0001100011100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100011100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001100011100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100011100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001100011100100) && ({row_reg, col_reg}<16'b0001100011100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100011100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100011100111) && ({row_reg, col_reg}<16'b0001100011101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100011101101) && ({row_reg, col_reg}<16'b0001100011110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001100011110000) && ({row_reg, col_reg}<16'b0001100011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100011110010) && ({row_reg, col_reg}<16'b0001100011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001100011111001) && ({row_reg, col_reg}<16'b0001100011111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0001100011111011) && ({row_reg, col_reg}<16'b0001100100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100100000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100100000001) && ({row_reg, col_reg}<16'b0001100100000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001100100000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001100100000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100100000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100100000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100100000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001100100001000) && ({row_reg, col_reg}<16'b0001100100001010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001100100001010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001100100001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001100100001100) && ({row_reg, col_reg}<16'b0001100100001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100100001110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001100100001111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001100100010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100100010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001100100010010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0001100100010011)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0001100100010100) && ({row_reg, col_reg}<16'b0001100100010110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0001100100010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100100010111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001100100011000) && ({row_reg, col_reg}<16'b0001100100011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100100011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001100100011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100100011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100100011101) && ({row_reg, col_reg}<16'b0001100100100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100100100000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001100100100001) && ({row_reg, col_reg}<16'b0001100100100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001100100100011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001100100100100) && ({row_reg, col_reg}<16'b0001100100100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100100100110)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0001100100100111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0001100100101000) && ({row_reg, col_reg}<16'b0001100100101010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001100100101010) && ({row_reg, col_reg}<16'b0001100100101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100100101101) && ({row_reg, col_reg}<16'b0001100100101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001100100101111) && ({row_reg, col_reg}<16'b0001100100110001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001100100110001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001100100110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100100110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001100100110100) && ({row_reg, col_reg}<16'b0001100100110110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001100100110110) && ({row_reg, col_reg}<16'b0001100100111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100100111001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001100100111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001100100111011) && ({row_reg, col_reg}<16'b0001100100111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100100111101) && ({row_reg, col_reg}<16'b0001100100111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100100111111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001100101000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001100101000001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0001100101000010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001100101000011) && ({row_reg, col_reg}<16'b0001100101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100101000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001100101000111) && ({row_reg, col_reg}<16'b0001100101001001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001100101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001100101001010) && ({row_reg, col_reg}<16'b0001100101001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100101001110) && ({row_reg, col_reg}<16'b0001100101010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100101010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001100101010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100101010010)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0001100101010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001100101010100) && ({row_reg, col_reg}<16'b0001100101010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100101010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100101010111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001100101011000) && ({row_reg, col_reg}<16'b0001100101011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100101011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001100101011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001100101011100) && ({row_reg, col_reg}<16'b0001100101011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100101011110) && ({row_reg, col_reg}<16'b0001100101100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100101100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001100101100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001100101100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001100101100110) && ({row_reg, col_reg}<16'b0001100101101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001100101101000) && ({row_reg, col_reg}<16'b0001100101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100101101010) && ({row_reg, col_reg}<16'b0001100101101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100101101101) && ({row_reg, col_reg}<16'b0001100101110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001100101110000) && ({row_reg, col_reg}<16'b0001100101110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100101110100) && ({row_reg, col_reg}<16'b0001100101111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100101111000) && ({row_reg, col_reg}<16'b0001100101111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100101111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100101111011) && ({row_reg, col_reg}<16'b0001100101111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100101111101) && ({row_reg, col_reg}<16'b0001100110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100110000010) && ({row_reg, col_reg}<16'b0001100110100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001100110100011) && ({row_reg, col_reg}<16'b0001100110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100110101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100110101011) && ({row_reg, col_reg}<16'b0001100110101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001100110101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001100110101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100110110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100110110001) && ({row_reg, col_reg}<16'b0001100110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001100110110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100110110100) && ({row_reg, col_reg}<16'b0001100110110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100110110111) && ({row_reg, col_reg}<16'b0001100110111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001100110111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100110111010) && ({row_reg, col_reg}<16'b0001100110111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100110111100) && ({row_reg, col_reg}<16'b0001100110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001100110111111) && ({row_reg, col_reg}<16'b0001100111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100111000101) && ({row_reg, col_reg}<16'b0001100111000111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001100111000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100111001000) && ({row_reg, col_reg}<16'b0001100111001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001100111001010) && ({row_reg, col_reg}<16'b0001100111001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001100111001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100111001110) && ({row_reg, col_reg}<16'b0001100111010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001100111010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100111010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001100111010101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001100111010110) && ({row_reg, col_reg}<16'b0001100111011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100111011000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0001100111011001) && ({row_reg, col_reg}<16'b0001100111011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100111011100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001100111011101) && ({row_reg, col_reg}<16'b0001100111100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100111100000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001100111100001) && ({row_reg, col_reg}<16'b0001100111100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100111100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001100111100100) && ({row_reg, col_reg}<16'b0001100111101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100111101101) && ({row_reg, col_reg}<16'b0001100111110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001100111110000) && ({row_reg, col_reg}<16'b0001100111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100111110010) && ({row_reg, col_reg}<16'b0001100111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001100111111001) && ({row_reg, col_reg}<16'b0001100111111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0001100111111011) && ({row_reg, col_reg}<16'b0001101000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101000000000) && ({row_reg, col_reg}<16'b0001101000000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101000000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101000000110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001101000000111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001101000001000) && ({row_reg, col_reg}<16'b0001101000001010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001101000001010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001101000001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101000001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001101000001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001101000001110) && ({row_reg, col_reg}<16'b0001101000010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101000010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001101000010001)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0001101000010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001101000010011)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0001101000010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101000010101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001101000010110) && ({row_reg, col_reg}<16'b0001101000011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101000011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001101000011001) && ({row_reg, col_reg}<16'b0001101000011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101000011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101000011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001101000011101) && ({row_reg, col_reg}<16'b0001101000011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101000011111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001101000100000) && ({row_reg, col_reg}<16'b0001101000100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001101000100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001101000100110) && ({row_reg, col_reg}<16'b0001101000101001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001101000101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101000101010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001101000101011) && ({row_reg, col_reg}<16'b0001101000101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101000101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001101000101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001101000101111) && ({row_reg, col_reg}<16'b0001101000110001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001101000110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101000110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001101000110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001101000110100) && ({row_reg, col_reg}<16'b0001101000110110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001101000110110) && ({row_reg, col_reg}<16'b0001101000111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101000111001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001101000111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001101000111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101000111100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101000111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101000111110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001101000111111) && ({row_reg, col_reg}<16'b0001101001000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001101001000001) && ({row_reg, col_reg}<16'b0001101001000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001101001000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101001000100)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}==16'b0001101001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101001000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001101001000111) && ({row_reg, col_reg}<16'b0001101001001001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001101001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001101001001100) && ({row_reg, col_reg}<16'b0001101001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101001010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0001101001010001) && ({row_reg, col_reg}<16'b0001101001010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001101001010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001101001010100) && ({row_reg, col_reg}<16'b0001101001010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101001010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001101001010111) && ({row_reg, col_reg}<16'b0001101001011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001101001011010) && ({row_reg, col_reg}<16'b0001101001011101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001101001011101) && ({row_reg, col_reg}<16'b0001101001011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101001100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001101001100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101001100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101001100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001101001100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101001100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001101001100110) && ({row_reg, col_reg}<16'b0001101001101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101001101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001101001101001) && ({row_reg, col_reg}<16'b0001101001101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001101001101011) && ({row_reg, col_reg}<16'b0001101001101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101001101101) && ({row_reg, col_reg}<16'b0001101001110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001101001110000) && ({row_reg, col_reg}<16'b0001101001110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101001110100) && ({row_reg, col_reg}<16'b0001101001110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001101001110110) && ({row_reg, col_reg}<16'b0001101001111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101001111000) && ({row_reg, col_reg}<16'b0001101001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101001111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101001111100) && ({row_reg, col_reg}<16'b0001101010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101010000010) && ({row_reg, col_reg}<16'b0001101010100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001101010100011) && ({row_reg, col_reg}<16'b0001101010100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101010100111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101010101000) && ({row_reg, col_reg}<16'b0001101010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101010101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001101010101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001101010101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001101010101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001101010101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001101010101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101010110000) && ({row_reg, col_reg}<16'b0001101010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001101010110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101010110100) && ({row_reg, col_reg}<16'b0001101010110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101010110111) && ({row_reg, col_reg}<16'b0001101010111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001101010111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101010111010) && ({row_reg, col_reg}<16'b0001101010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101010111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001101010111101) && ({row_reg, col_reg}<16'b0001101011000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001101011000000) && ({row_reg, col_reg}<16'b0001101011000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101011000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001101011000110) && ({row_reg, col_reg}<16'b0001101011001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001101011001000) && ({row_reg, col_reg}<16'b0001101011001100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001101011001100) && ({row_reg, col_reg}<16'b0001101011010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001101011010101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001101011010110) && ({row_reg, col_reg}<16'b0001101011011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101011011000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0001101011011001) && ({row_reg, col_reg}<16'b0001101011011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101011011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001101011011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001101011011101) && ({row_reg, col_reg}<16'b0001101011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101011011111) && ({row_reg, col_reg}<16'b0001101011100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001101011100001) && ({row_reg, col_reg}<16'b0001101011100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101011100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001101011100100) && ({row_reg, col_reg}<16'b0001101011101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101011101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001101011101001) && ({row_reg, col_reg}<16'b0001101011101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001101011101101) && ({row_reg, col_reg}<16'b0001101011110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001101011110000) && ({row_reg, col_reg}<16'b0001101011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101011110010) && ({row_reg, col_reg}<16'b0001101011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001101011111001) && ({row_reg, col_reg}<16'b0001101011111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0001101011111011) && ({row_reg, col_reg}<16'b0001101100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101100000000) && ({row_reg, col_reg}<16'b0001101100000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101100000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101100000110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001101100000111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001101100001000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0001101100001001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001101100001010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001101100001011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001101100001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101100001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001101100001110) && ({row_reg, col_reg}<16'b0001101100010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101100010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001101100010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001101100010010) && ({row_reg, col_reg}<16'b0001101100010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001101100010100) && ({row_reg, col_reg}<16'b0001101100011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101100011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001101100011001) && ({row_reg, col_reg}<16'b0001101100011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101100011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101100011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001101100011101) && ({row_reg, col_reg}<16'b0001101100100000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001101100100000) && ({row_reg, col_reg}<16'b0001101100100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001101100100101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001101100100110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001101100100111)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0001101100101000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001101100101001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001101100101010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101100101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101100101100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001101100101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001101100101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001101100101111) && ({row_reg, col_reg}<16'b0001101100110001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001101100110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101100110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101100110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001101100110100) && ({row_reg, col_reg}<16'b0001101100110110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001101100110110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001101100110111) && ({row_reg, col_reg}<16'b0001101100111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101100111010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0001101100111011) && ({row_reg, col_reg}<16'b0001101100111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101100111101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001101100111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101100111111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001101101000000) && ({row_reg, col_reg}<16'b0001101101000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001101101000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101101000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101101000111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001101101001000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001101101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101101001010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001101101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001101101001100) && ({row_reg, col_reg}<16'b0001101101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101101010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001101101010001) && ({row_reg, col_reg}<16'b0001101101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001101101010100) && ({row_reg, col_reg}<16'b0001101101010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101101010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001101101010111) && ({row_reg, col_reg}<16'b0001101101011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001101101011010) && ({row_reg, col_reg}<16'b0001101101011100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001101101011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101101011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001101101011110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001101101011111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0001101101100000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001101101100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001101101100010) && ({row_reg, col_reg}<16'b0001101101100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101101100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101101100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001101101100110) && ({row_reg, col_reg}<16'b0001101101101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001101101101001) && ({row_reg, col_reg}<16'b0001101101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101101101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101101101101) && ({row_reg, col_reg}<16'b0001101101110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001101101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101101110001) && ({row_reg, col_reg}<16'b0001101101111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101101111000) && ({row_reg, col_reg}<16'b0001101101111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101101111010) && ({row_reg, col_reg}<16'b0001101101111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101101111100) && ({row_reg, col_reg}<16'b0001101110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101110000010) && ({row_reg, col_reg}<16'b0001101110100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001101110100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101110100100) && ({row_reg, col_reg}<16'b0001101110100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101110100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001101110101000) && ({row_reg, col_reg}<16'b0001101110101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001101110101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001101110101011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=16'b0001101110101100) && ({row_reg, col_reg}<16'b0001101110101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101110101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001101110101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101110110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101110110001) && ({row_reg, col_reg}<16'b0001101110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001101110110011) && ({row_reg, col_reg}<16'b0001101110110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101110110111) && ({row_reg, col_reg}<16'b0001101110111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001101110111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101110111010) && ({row_reg, col_reg}<16'b0001101110111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001101110111100) && ({row_reg, col_reg}<16'b0001101110111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001101110111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001101110111111) && ({row_reg, col_reg}<16'b0001101111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101111000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001101111000110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0001101111000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001101111001000) && ({row_reg, col_reg}<16'b0001101111001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001101111001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001101111001011) && ({row_reg, col_reg}<16'b0001101111001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001101111001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101111001110) && ({row_reg, col_reg}<16'b0001101111010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001101111010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101111010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001101111010110) && ({row_reg, col_reg}<16'b0001101111011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001101111011010) && ({row_reg, col_reg}<16'b0001101111011100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001101111011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001101111011101) && ({row_reg, col_reg}<16'b0001101111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101111011111) && ({row_reg, col_reg}<16'b0001101111100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001101111100001) && ({row_reg, col_reg}<16'b0001101111100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101111100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001101111100100) && ({row_reg, col_reg}<16'b0001101111101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001101111101101) && ({row_reg, col_reg}<16'b0001101111110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001101111110000) && ({row_reg, col_reg}<16'b0001101111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101111110010) && ({row_reg, col_reg}<16'b0001101111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001101111111001) && ({row_reg, col_reg}<16'b0001101111111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0001101111111011) && ({row_reg, col_reg}<16'b0001110000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110000000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001110000000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001110000000010) && ({row_reg, col_reg}<16'b0001110000000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110000000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110000000110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001110000000111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001110000001000) && ({row_reg, col_reg}<16'b0001110000001011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001110000001011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001110000001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110000001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001110000001110) && ({row_reg, col_reg}<16'b0001110000010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110000010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110000010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110000010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001110000010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001110000010100) && ({row_reg, col_reg}<16'b0001110000010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110000010111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001110000011000) && ({row_reg, col_reg}<16'b0001110000011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110000011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001110000011100) && ({row_reg, col_reg}<16'b0001110000011110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001110000011110) && ({row_reg, col_reg}<16'b0001110000100000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001110000100000) && ({row_reg, col_reg}<16'b0001110000100010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0001110000100010)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0001110000100011) && ({row_reg, col_reg}<16'b0001110000100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001110000100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001110000100110) && ({row_reg, col_reg}<16'b0001110000101001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001110000101001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001110000101010) && ({row_reg, col_reg}<16'b0001110000101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110000101100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001110000101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001110000101110) && ({row_reg, col_reg}<16'b0001110000110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001110000110001) && ({row_reg, col_reg}<16'b0001110000110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110000110011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001110000110100) && ({row_reg, col_reg}<16'b0001110000110110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001110000110110) && ({row_reg, col_reg}<16'b0001110000111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110000111010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001110000111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001110000111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110000111101) && ({row_reg, col_reg}<16'b0001110001000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001110001000000) && ({row_reg, col_reg}<16'b0001110001000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001110001000011) && ({row_reg, col_reg}<16'b0001110001000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110001000110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001110001000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110001001000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001110001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110001001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001110001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110001001100) && ({row_reg, col_reg}<16'b0001110001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110001010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0001110001010001) && ({row_reg, col_reg}<16'b0001110001010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001110001010011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0001110001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001110001010101) && ({row_reg, col_reg}<16'b0001110001010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110001010111) && ({row_reg, col_reg}<16'b0001110001011001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001110001011001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001110001011010) && ({row_reg, col_reg}<16'b0001110001011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110001011100) && ({row_reg, col_reg}<16'b0001110001011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001110001011110) && ({row_reg, col_reg}<16'b0001110001100000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001110001100000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0001110001100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110001100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110001100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001110001100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110001100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001110001100110) && ({row_reg, col_reg}<16'b0001110001101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110001101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001110001101001) && ({row_reg, col_reg}<16'b0001110001101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110001101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110001101101) && ({row_reg, col_reg}<16'b0001110001110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001110001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110001110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110001110010) && ({row_reg, col_reg}<16'b0001110001110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001110001110100) && ({row_reg, col_reg}<16'b0001110001111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110001111000) && ({row_reg, col_reg}<16'b0001110001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110001111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110001111100) && ({row_reg, col_reg}<16'b0001110001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110010000000) && ({row_reg, col_reg}<16'b0001110010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110010000011) && ({row_reg, col_reg}<16'b0001110010100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001110010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110010100101) && ({row_reg, col_reg}<16'b0001110010100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110010100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001110010101000) && ({row_reg, col_reg}<16'b0001110010101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001110010101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001110010101100) && ({row_reg, col_reg}<16'b0001110010101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001110010101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110010110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110010110001) && ({row_reg, col_reg}<16'b0001110010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001110010110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110010110100) && ({row_reg, col_reg}<16'b0001110010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001110010110110) && ({row_reg, col_reg}<16'b0001110010111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110010111000) && ({row_reg, col_reg}<16'b0001110010111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001110010111010) && ({row_reg, col_reg}<16'b0001110010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001110010111101) && ({row_reg, col_reg}<16'b0001110010111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001110011000000) && ({row_reg, col_reg}<16'b0001110011000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110011000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001110011000110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0001110011000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110011001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001110011001001) && ({row_reg, col_reg}<16'b0001110011001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110011001011) && ({row_reg, col_reg}<16'b0001110011001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001110011001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110011001110) && ({row_reg, col_reg}<16'b0001110011010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001110011010100) && ({row_reg, col_reg}<16'b0001110011010110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001110011010110) && ({row_reg, col_reg}<16'b0001110011011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001110011011000) && ({row_reg, col_reg}<16'b0001110011011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110011011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110011011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001110011011101) && ({row_reg, col_reg}<16'b0001110011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110011011111) && ({row_reg, col_reg}<16'b0001110011100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001110011100001) && ({row_reg, col_reg}<16'b0001110011100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110011100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001110011100100) && ({row_reg, col_reg}<16'b0001110011101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110011101101) && ({row_reg, col_reg}<16'b0001110011110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001110011110000) && ({row_reg, col_reg}<16'b0001110011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110011110010) && ({row_reg, col_reg}<16'b0001110011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001110011111001) && ({row_reg, col_reg}<16'b0001110011111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0001110011111011) && ({row_reg, col_reg}<16'b0001110100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110100000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001110100000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001110100000010) && ({row_reg, col_reg}<16'b0001110100000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110100000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110100000110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001110100000111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001110100001000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001110100001001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0001110100001010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001110100001011) && ({row_reg, col_reg}<16'b0001110100001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110100001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001110100001110) && ({row_reg, col_reg}<16'b0001110100010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001110100010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110100010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110100010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001110100010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001110100010100) && ({row_reg, col_reg}<16'b0001110100010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110100010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001110100010111) && ({row_reg, col_reg}<16'b0001110100011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110100011001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001110100011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001110100011011) && ({row_reg, col_reg}<16'b0001110100011111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001110100011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001110100100000) && ({row_reg, col_reg}<16'b0001110100100010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0001110100100010)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0001110100100011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0001110100100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001110100100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110100100110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001110100100111) && ({row_reg, col_reg}<16'b0001110100101001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001110100101001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001110100101010) && ({row_reg, col_reg}<16'b0001110100101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110100101100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001110100101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001110100101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110100101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001110100110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110100110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110100110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110100110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001110100110100) && ({row_reg, col_reg}<16'b0001110100111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110100111010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0001110100111011) && ({row_reg, col_reg}<16'b0001110100111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110100111101) && ({row_reg, col_reg}<16'b0001110101000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110101000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001110101000001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0001110101000010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001110101000011) && ({row_reg, col_reg}<16'b0001110101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110101000110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001110101000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110101001000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001110101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110101001010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0001110101001011) && ({row_reg, col_reg}<16'b0001110101001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110101001101) && ({row_reg, col_reg}<16'b0001110101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001110101010000) && ({row_reg, col_reg}<16'b0001110101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001110101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001110101010101) && ({row_reg, col_reg}<16'b0001110101010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110101010111) && ({row_reg, col_reg}<16'b0001110101011001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001110101011001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110101011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110101011011) && ({row_reg, col_reg}<16'b0001110101011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001110101011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110101011110) && ({row_reg, col_reg}<16'b0001110101100001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001110101100001)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0001110101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110101100011) && ({row_reg, col_reg}<16'b0001110101100110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110101100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110101100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001110101101000) && ({row_reg, col_reg}<16'b0001110101101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001110101101101) && ({row_reg, col_reg}<16'b0001110101110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001110101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110101110001) && ({row_reg, col_reg}<16'b0001110101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001110101110100) && ({row_reg, col_reg}<16'b0001110101111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110101111000) && ({row_reg, col_reg}<16'b0001110101111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110101111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110101111100) && ({row_reg, col_reg}<16'b0001110101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001110101111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001110110000000) && ({row_reg, col_reg}<16'b0001110110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110110000011) && ({row_reg, col_reg}<16'b0001110110100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001110110100100) && ({row_reg, col_reg}<16'b0001110110100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110110100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110110100111) && ({row_reg, col_reg}<16'b0001110110101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001110110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110110101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110110101100) && ({row_reg, col_reg}<16'b0001110110101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001110110101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001110110101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110110110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110110110001) && ({row_reg, col_reg}<16'b0001110110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001110110110011) && ({row_reg, col_reg}<16'b0001110110110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110110110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110110111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001110110111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110110111010) && ({row_reg, col_reg}<16'b0001110110111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001110110111110) && ({row_reg, col_reg}<16'b0001110111000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001110111000000) && ({row_reg, col_reg}<16'b0001110111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110111000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001110111000110) && ({row_reg, col_reg}<16'b0001110111001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110111001011) && ({row_reg, col_reg}<16'b0001110111001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001110111001101) && ({row_reg, col_reg}<16'b0001110111001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110111001111) && ({row_reg, col_reg}<16'b0001110111010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001110111010010) && ({row_reg, col_reg}<16'b0001110111010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110111010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110111010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110111010110) && ({row_reg, col_reg}<16'b0001110111011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001110111011000) && ({row_reg, col_reg}<16'b0001110111011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110111011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001110111011101) && ({row_reg, col_reg}<16'b0001110111100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110111100000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001110111100001) && ({row_reg, col_reg}<16'b0001110111100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110111100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001110111100100) && ({row_reg, col_reg}<16'b0001110111101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110111101101) && ({row_reg, col_reg}<16'b0001110111110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001110111110000) && ({row_reg, col_reg}<16'b0001110111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110111110010) && ({row_reg, col_reg}<16'b0001110111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001110111111001) && ({row_reg, col_reg}<16'b0001110111111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0001110111111011) && ({row_reg, col_reg}<16'b0001111000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111000000000)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}>=16'b0001111000000001) && ({row_reg, col_reg}<16'b0001111000000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001111000000100) && ({row_reg, col_reg}<16'b0001111000000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111000000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111000000111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001111000001000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001111000001001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001111000001010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001111000001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111000001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001111000001101) && ({row_reg, col_reg}<16'b0001111000010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111000010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111000010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001111000010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001111000010100) && ({row_reg, col_reg}<16'b0001111000010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111000010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001111000010111) && ({row_reg, col_reg}<16'b0001111000011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111000011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111000011010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001111000011011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001111000011100) && ({row_reg, col_reg}<16'b0001111000100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111000100000)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0001111000100001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0001111000100010) && ({row_reg, col_reg}<16'b0001111000100100)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0001111000100100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0001111000100101) && ({row_reg, col_reg}<16'b0001111000100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111000100111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001111000101000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001111000101001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001111000101010) && ({row_reg, col_reg}<16'b0001111000101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111000101100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001111000101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001111000101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111000101111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001111000110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111000110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111000110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111000110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111000110100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001111000110101) && ({row_reg, col_reg}<16'b0001111000110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001111000110111) && ({row_reg, col_reg}<16'b0001111000111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111000111001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001111000111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001111000111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001111000111100) && ({row_reg, col_reg}<16'b0001111000111110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111000111110) && ({row_reg, col_reg}<16'b0001111001000000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001111001000000) && ({row_reg, col_reg}<16'b0001111001000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001111001000011) && ({row_reg, col_reg}<16'b0001111001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111001000110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001111001000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111001001000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001111001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111001001010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001111001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001111001001100) && ({row_reg, col_reg}<16'b0001111001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111001010000) && ({row_reg, col_reg}<16'b0001111001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001111001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111001010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111001010110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0001111001010111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111001011000) && ({row_reg, col_reg}<16'b0001111001011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001111001011010) && ({row_reg, col_reg}<16'b0001111001011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001111001011100) && ({row_reg, col_reg}<16'b0001111001011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111001011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111001011111) && ({row_reg, col_reg}<16'b0001111001100010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001111001100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001111001100011) && ({row_reg, col_reg}<16'b0001111001100110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001111001100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111001100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001111001101000) && ({row_reg, col_reg}<16'b0001111001101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001111001101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111001101110) && ({row_reg, col_reg}<16'b0001111001110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111001110000) && ({row_reg, col_reg}<16'b0001111001110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111001110010) && ({row_reg, col_reg}<16'b0001111001110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001111001110100) && ({row_reg, col_reg}<16'b0001111001111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001111001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111001111001) && ({row_reg, col_reg}<16'b0001111001111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111001111100) && ({row_reg, col_reg}<16'b0001111001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001111001111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001111010000000) && ({row_reg, col_reg}<16'b0001111010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111010000011) && ({row_reg, col_reg}<16'b0001111010100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001111010100011) && ({row_reg, col_reg}<16'b0001111010100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001111010100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111010100111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111010101000) && ({row_reg, col_reg}<16'b0001111010101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111010101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111010101100) && ({row_reg, col_reg}<16'b0001111010101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001111010101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001111010101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111010110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111010110001) && ({row_reg, col_reg}<16'b0001111010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001111010110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111010110100) && ({row_reg, col_reg}<16'b0001111010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111010110110) && ({row_reg, col_reg}<16'b0001111010111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111010111010) && ({row_reg, col_reg}<16'b0001111010111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111010111110) && ({row_reg, col_reg}<16'b0001111011000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001111011000000) && ({row_reg, col_reg}<16'b0001111011000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111011000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111011000110) && ({row_reg, col_reg}<16'b0001111011001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111011001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111011001100) && ({row_reg, col_reg}<16'b0001111011010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111011010000) && ({row_reg, col_reg}<16'b0001111011010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001111011010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111011010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001111011010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001111011010110) && ({row_reg, col_reg}<16'b0001111011011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001111011011000) && ({row_reg, col_reg}<16'b0001111011011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111011011010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0001111011011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111011011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111011011101) && ({row_reg, col_reg}<16'b0001111011100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111011100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111011100100) && ({row_reg, col_reg}<16'b0001111011101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111011101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111011101001) && ({row_reg, col_reg}<16'b0001111011101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001111011101101) && ({row_reg, col_reg}<16'b0001111011110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111011110000) && ({row_reg, col_reg}<16'b0001111011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111011110010) && ({row_reg, col_reg}<16'b0001111011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001111011111001)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0001111011111010) && ({row_reg, col_reg}<16'b0001111100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111100000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001111100000001) && ({row_reg, col_reg}<16'b0001111100000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111100000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001111100000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111100000111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001111100001000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001111100001001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001111100001010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001111100001011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001111100001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001111100001101) && ({row_reg, col_reg}<16'b0001111100001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111100001111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001111100010000) && ({row_reg, col_reg}<16'b0001111100010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111100010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001111100010011) && ({row_reg, col_reg}<16'b0001111100010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001111100010101) && ({row_reg, col_reg}<16'b0001111100010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001111100010111) && ({row_reg, col_reg}<16'b0001111100011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111100011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111100011010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001111100011011)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0001111100011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001111100011101) && ({row_reg, col_reg}<16'b0001111100100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001111100100000) && ({row_reg, col_reg}<16'b0001111100100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001111100100101) && ({row_reg, col_reg}<16'b0001111100100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111100100111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001111100101000) && ({row_reg, col_reg}<16'b0001111100101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001111100101010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001111100101011) && ({row_reg, col_reg}<16'b0001111100101110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001111100101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111100101111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001111100110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111100110001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001111100110010) && ({row_reg, col_reg}<16'b0001111100110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111100110100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001111100110101) && ({row_reg, col_reg}<16'b0001111100110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001111100110111) && ({row_reg, col_reg}<16'b0001111100111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001111100111001) && ({row_reg, col_reg}<16'b0001111100111011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001111100111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001111100111100) && ({row_reg, col_reg}<16'b0001111100111110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111100111110) && ({row_reg, col_reg}<16'b0001111101000000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001111101000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001111101000001) && ({row_reg, col_reg}<16'b0001111101000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001111101000011) && ({row_reg, col_reg}<16'b0001111101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111101000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111101000111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001111101001000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001111101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001111101001100) && ({row_reg, col_reg}<16'b0001111101010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111101010001) && ({row_reg, col_reg}<16'b0001111101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001111101010100) && ({row_reg, col_reg}<16'b0001111101010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111101010110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0001111101010111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001111101011000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001111101011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111101011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001111101011011) && ({row_reg, col_reg}<16'b0001111101011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111101011111) && ({row_reg, col_reg}<16'b0001111101100010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001111101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111101100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111101100100) && ({row_reg, col_reg}<16'b0001111101100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111101100110) && ({row_reg, col_reg}<16'b0001111101101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001111101101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001111101101001) && ({row_reg, col_reg}<16'b0001111101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111101101110) && ({row_reg, col_reg}<16'b0001111101110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111101110000) && ({row_reg, col_reg}<16'b0001111101110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111101110010) && ({row_reg, col_reg}<16'b0001111101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001111101110100) && ({row_reg, col_reg}<16'b0001111101111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001111101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111101111001) && ({row_reg, col_reg}<16'b0001111101111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111101111100) && ({row_reg, col_reg}<16'b0001111101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111101111110) && ({row_reg, col_reg}<16'b0001111110000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001111110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001111110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111110000011) && ({row_reg, col_reg}<16'b0001111110100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001111110100011) && ({row_reg, col_reg}<16'b0001111110100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001111110100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111110100111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111110101000) && ({row_reg, col_reg}<16'b0001111110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111110101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111110101100) && ({row_reg, col_reg}<16'b0001111110101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001111110101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001111110101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111110110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111110110001) && ({row_reg, col_reg}<16'b0001111110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001111110110011) && ({row_reg, col_reg}<16'b0001111110111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111110111010) && ({row_reg, col_reg}<16'b0001111110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111110111101) && ({row_reg, col_reg}<16'b0001111111000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001111111000000) && ({row_reg, col_reg}<16'b0001111111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111111000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111111000110) && ({row_reg, col_reg}<16'b0001111111001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111111001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111111001100) && ({row_reg, col_reg}<16'b0001111111010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111111010000) && ({row_reg, col_reg}<16'b0001111111010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111111010101) && ({row_reg, col_reg}<16'b0001111111011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111111011010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0001111111011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111111011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111111011101) && ({row_reg, col_reg}<16'b0001111111100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111111100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111111100100) && ({row_reg, col_reg}<16'b0001111111101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111111101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111111101001) && ({row_reg, col_reg}<16'b0001111111101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001111111101101) && ({row_reg, col_reg}<16'b0001111111101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111111101111) && ({row_reg, col_reg}<16'b0001111111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111111110010) && ({row_reg, col_reg}<16'b0001111111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001111111111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111111111010) && ({row_reg, col_reg}<16'b0001111111111111)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}==16'b0001111111111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000000000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010000000000001) && ({row_reg, col_reg}<16'b0010000000000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000000000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010000000000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000000000111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010000000001000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0010000000001001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010000000001010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0010000000001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000000001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0010000000001101) && ({row_reg, col_reg}<16'b0010000000010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000000010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010000000010011) && ({row_reg, col_reg}<16'b0010000000010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010000000010101) && ({row_reg, col_reg}<16'b0010000000010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010000000010111) && ({row_reg, col_reg}<16'b0010000000011001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010000000011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000000011010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010000000011011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010000000011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010000000011101) && ({row_reg, col_reg}<16'b0010000000011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000000011111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010000000100000) && ({row_reg, col_reg}<16'b0010000000100010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010000000100010)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0010000000100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010000000100100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010000000100101) && ({row_reg, col_reg}<16'b0010000000100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010000000100111) && ({row_reg, col_reg}<16'b0010000000101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010000000101010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010000000101011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010000000101100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010000000101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010000000101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000000101111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010000000110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010000000110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000000110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000000110011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010000000110100) && ({row_reg, col_reg}<16'b0010000000110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000000110110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010000000110111) && ({row_reg, col_reg}<16'b0010000000111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000000111010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010000000111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010000000111100) && ({row_reg, col_reg}<16'b0010000000111110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000000111110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010000000111111) && ({row_reg, col_reg}<16'b0010000001000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000001000001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010000001000010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010000001000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010000001000100) && ({row_reg, col_reg}<16'b0010000001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000001000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010000001000111) && ({row_reg, col_reg}<16'b0010000001001001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010000001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010000001001100) && ({row_reg, col_reg}<16'b0010000001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000001010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000001010001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010000001010010) && ({row_reg, col_reg}<16'b0010000001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010000001010100) && ({row_reg, col_reg}<16'b0010000001010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000001010110) && ({row_reg, col_reg}<16'b0010000001011000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0010000001011000) && ({row_reg, col_reg}<16'b0010000001011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010000001011100) && ({row_reg, col_reg}<16'b0010000001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000001011111) && ({row_reg, col_reg}<16'b0010000001100010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010000001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000001100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000001100100) && ({row_reg, col_reg}<16'b0010000001100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000001100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010000001101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000001101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010000001101010) && ({row_reg, col_reg}<16'b0010000001101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010000001101110) && ({row_reg, col_reg}<16'b0010000001110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000001110000) && ({row_reg, col_reg}<16'b0010000001110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000001110010) && ({row_reg, col_reg}<16'b0010000001111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000001111000) && ({row_reg, col_reg}<16'b0010000001111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000001111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000001111100) && ({row_reg, col_reg}<16'b0010000001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000001111110) && ({row_reg, col_reg}<16'b0010000010000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010000010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010000010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000010000011) && ({row_reg, col_reg}<16'b0010000010100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010000010100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000010100100) && ({row_reg, col_reg}<16'b0010000010100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000010100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000010100111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000010101000) && ({row_reg, col_reg}<16'b0010000010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000010101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000010101110) && ({row_reg, col_reg}<16'b0010000010110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000010110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000010110001) && ({row_reg, col_reg}<16'b0010000010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010000010110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000010110100) && ({row_reg, col_reg}<16'b0010000010111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000010111010) && ({row_reg, col_reg}<16'b0010000010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010000010111101) && ({row_reg, col_reg}<16'b0010000010111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010000010111111) && ({row_reg, col_reg}<16'b0010000011000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000011000001) && ({row_reg, col_reg}<16'b0010000011000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000011000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000011000110) && ({row_reg, col_reg}<16'b0010000011001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000011001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000011001100) && ({row_reg, col_reg}<16'b0010000011010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000011010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010000011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000011010010) && ({row_reg, col_reg}<16'b0010000011010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010000011010101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010000011010110) && ({row_reg, col_reg}<16'b0010000011011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000011011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000011011101) && ({row_reg, col_reg}<16'b0010000011100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000011100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010000011100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000011100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000011100100) && ({row_reg, col_reg}<16'b0010000011101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000011101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000011101110) && ({row_reg, col_reg}<16'b0010000011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000011110010) && ({row_reg, col_reg}<16'b0010000011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010000011111001) && ({row_reg, col_reg}<16'b0010000011111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000011111011) && ({row_reg, col_reg}<16'b0010000011111110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0010000011111110) && ({row_reg, col_reg}<16'b0010000100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000100000000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010000100000001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010000100000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000100000011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010000100000100) && ({row_reg, col_reg}<16'b0010000100000110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010000100000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000100000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010000100001000) && ({row_reg, col_reg}<16'b0010000100001010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010000100001010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010000100001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000100001100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010000100001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000100001110) && ({row_reg, col_reg}<16'b0010000100010000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010000100010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000100010001) && ({row_reg, col_reg}<16'b0010000100010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000100010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010000100010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010000100010101) && ({row_reg, col_reg}<16'b0010000100010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000100010111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010000100011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000100011001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010000100011010) && ({row_reg, col_reg}<16'b0010000100011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010000100011100) && ({row_reg, col_reg}<16'b0010000100011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010000100011110) && ({row_reg, col_reg}<16'b0010000100100000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010000100100000) && ({row_reg, col_reg}<16'b0010000100100010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010000100100010)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0010000100100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010000100100100) && ({row_reg, col_reg}<16'b0010000100100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000100100110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010000100100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010000100101000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0010000100101001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0010000100101010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010000100101011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010000100101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000100101101)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010000100101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010000100101111) && ({row_reg, col_reg}<16'b0010000100110001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010000100110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010000100110010) && ({row_reg, col_reg}<16'b0010000100110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000100110100) && ({row_reg, col_reg}<16'b0010000100110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000100110111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0010000100111000) && ({row_reg, col_reg}<16'b0010000100111010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010000100111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000100111011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010000100111100) && ({row_reg, col_reg}<16'b0010000100111110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010000100111110) && ({row_reg, col_reg}<16'b0010000101000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000101000001) && ({row_reg, col_reg}<16'b0010000101000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010000101000011) && ({row_reg, col_reg}<16'b0010000101000101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010000101000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010000101000110) && ({row_reg, col_reg}<16'b0010000101001000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000101001000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010000101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000101001010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010000101001011) && ({row_reg, col_reg}<16'b0010000101001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000101001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000101001110) && ({row_reg, col_reg}<16'b0010000101010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000101010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010000101010001) && ({row_reg, col_reg}<16'b0010000101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010000101010100) && ({row_reg, col_reg}<16'b0010000101010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000101010110) && ({row_reg, col_reg}<16'b0010000101011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010000101011011) && ({row_reg, col_reg}<16'b0010000101100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000101100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000101100001)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010000101100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000101100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010000101100100) && ({row_reg, col_reg}<16'b0010000101100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000101100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010000101101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000101101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010000101101010) && ({row_reg, col_reg}<16'b0010000101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010000101101110) && ({row_reg, col_reg}<16'b0010000101110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000101110000) && ({row_reg, col_reg}<16'b0010000101110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000101110010) && ({row_reg, col_reg}<16'b0010000101111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010000101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000101111001) && ({row_reg, col_reg}<16'b0010000101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000101111100) && ({row_reg, col_reg}<16'b0010000101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000101111110) && ({row_reg, col_reg}<16'b0010000110000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010000110000000) && ({row_reg, col_reg}<16'b0010000110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000110000011) && ({row_reg, col_reg}<16'b0010000110100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010000110100100) && ({row_reg, col_reg}<16'b0010000110100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000110100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000110100111) && ({row_reg, col_reg}<16'b0010000110101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000110101011) && ({row_reg, col_reg}<16'b0010000110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010000110110000) && ({row_reg, col_reg}<16'b0010000110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010000110110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000110110100) && ({row_reg, col_reg}<16'b0010000110111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000110111010) && ({row_reg, col_reg}<16'b0010000110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000110111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010000110111110) && ({row_reg, col_reg}<16'b0010000111000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000111000001) && ({row_reg, col_reg}<16'b0010000111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000111000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000111000110) && ({row_reg, col_reg}<16'b0010000111001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000111001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000111001100) && ({row_reg, col_reg}<16'b0010000111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000111001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010000111001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000111010000) && ({row_reg, col_reg}<16'b0010000111010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000111010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000111010011) && ({row_reg, col_reg}<16'b0010000111010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010000111010101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010000111010110) && ({row_reg, col_reg}<16'b0010000111011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010000111011011) && ({row_reg, col_reg}<16'b0010000111011101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010000111011101) && ({row_reg, col_reg}<16'b0010000111100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000111100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010000111100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000111100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000111100100) && ({row_reg, col_reg}<16'b0010000111101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000111101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000111101110) && ({row_reg, col_reg}<16'b0010000111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000111110010) && ({row_reg, col_reg}<16'b0010000111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010000111111001) && ({row_reg, col_reg}<16'b0010000111111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000111111011) && ({row_reg, col_reg}<16'b0010000111111110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0010000111111110) && ({row_reg, col_reg}<16'b0010001000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001000000000) && ({row_reg, col_reg}<16'b0010001000000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010001000000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001000000011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010001000000100)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0010001000000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001000000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001000000111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010001000001000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0010001000001001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010001000001010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010001000001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001000001100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010001000001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010001000001110) && ({row_reg, col_reg}<16'b0010001000010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001000010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001000010001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010001000010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001000010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010001000010100) && ({row_reg, col_reg}<16'b0010001000010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001000010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001000010111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010001000011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001000011001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010001000011010) && ({row_reg, col_reg}<16'b0010001000011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010001000011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010001000011101) && ({row_reg, col_reg}<16'b0010001000011111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010001000011111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010001000100000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010001000100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010001000100010) && ({row_reg, col_reg}<16'b0010001000100100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0010001000100100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010001000100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001000100110)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0010001000100111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0010001000101000) && ({row_reg, col_reg}<16'b0010001000101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010001000101010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010001000101011) && ({row_reg, col_reg}<16'b0010001000101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001000101101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010001000101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010001000101111) && ({row_reg, col_reg}<16'b0010001000110001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010001000110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010001000110010) && ({row_reg, col_reg}<16'b0010001000110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010001000110100) && ({row_reg, col_reg}<16'b0010001000111000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010001000111000) && ({row_reg, col_reg}<16'b0010001000111100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010001000111100) && ({row_reg, col_reg}<16'b0010001000111111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001000111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001001000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010001001000001) && ({row_reg, col_reg}<16'b0010001001000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001001000011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010001001000100) && ({row_reg, col_reg}<16'b0010001001000110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010001001000110) && ({row_reg, col_reg}<16'b0010001001001000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001001001000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010001001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001001001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010001001001011) && ({row_reg, col_reg}<16'b0010001001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001001001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010001001010000) && ({row_reg, col_reg}<16'b0010001001010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001001010010)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0010001001010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010001001010101) && ({row_reg, col_reg}<16'b0010001001011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001001011000) && ({row_reg, col_reg}<16'b0010001001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001001011111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010001001100000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010001001100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010001001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001001100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010001001100100) && ({row_reg, col_reg}<16'b0010001001100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010001001100110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010001001100111) && ({row_reg, col_reg}<16'b0010001001101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001001101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010001001101010) && ({row_reg, col_reg}<16'b0010001001101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010001001101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010001001101110) && ({row_reg, col_reg}<16'b0010001001110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001001110000) && ({row_reg, col_reg}<16'b0010001001110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001001110010) && ({row_reg, col_reg}<16'b0010001001110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010001001110100) && ({row_reg, col_reg}<16'b0010001001110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001001110111) && ({row_reg, col_reg}<16'b0010001001111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001001111001) && ({row_reg, col_reg}<16'b0010001001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010001001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001001111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010001001111101) && ({row_reg, col_reg}<16'b0010001010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001010000000) && ({row_reg, col_reg}<16'b0010001010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001010000011) && ({row_reg, col_reg}<16'b0010001010100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010001010100100) && ({row_reg, col_reg}<16'b0010001010101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001010101000) && ({row_reg, col_reg}<16'b0010001010101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001010101011) && ({row_reg, col_reg}<16'b0010001010101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010001010101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001010110000) && ({row_reg, col_reg}<16'b0010001010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010001010110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001010110100) && ({row_reg, col_reg}<16'b0010001010111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001010111010) && ({row_reg, col_reg}<16'b0010001010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001010111101) && ({row_reg, col_reg}<16'b0010001010111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010001010111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001011000000) && ({row_reg, col_reg}<16'b0010001011000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001011000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001011000110) && ({row_reg, col_reg}<16'b0010001011001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001011001011) && ({row_reg, col_reg}<16'b0010001011001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010001011001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001011001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001011001111) && ({row_reg, col_reg}<16'b0010001011010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010001011010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001011010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010001011010101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010001011010110) && ({row_reg, col_reg}<16'b0010001011011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001011011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010001011011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001011011101) && ({row_reg, col_reg}<16'b0010001011100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001011100000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001011100001) && ({row_reg, col_reg}<16'b0010001011100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001011100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001011100100) && ({row_reg, col_reg}<16'b0010001011101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001011101010) && ({row_reg, col_reg}<16'b0010001011101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001011101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001011101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001011101110) && ({row_reg, col_reg}<16'b0010001011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001011110010) && ({row_reg, col_reg}<16'b0010001011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010001011111001) && ({row_reg, col_reg}<16'b0010001011111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001011111011) && ({row_reg, col_reg}<16'b0010001011111111)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}==16'b0010001011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001100000000) && ({row_reg, col_reg}<16'b0010001100000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010001100000010) && ({row_reg, col_reg}<16'b0010001100000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001100000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010001100000110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001100000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010001100001000) && ({row_reg, col_reg}<16'b0010001100001011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010001100001011) && ({row_reg, col_reg}<16'b0010001100010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001100010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001100010011) && ({row_reg, col_reg}<16'b0010001100010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010001100010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001100010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010001100010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001100011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001100011001)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0010001100011010) && ({row_reg, col_reg}<16'b0010001100011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010001100011100) && ({row_reg, col_reg}<16'b0010001100011110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010001100011110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010001100011111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010001100100000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010001100100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010001100100010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0010001100100011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010001100100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010001100100101) && ({row_reg, col_reg}<16'b0010001100100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001100100111)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0010001100101000)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0010001100101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001100101010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001100101011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010001100101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001100101101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010001100101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001100101111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010001100110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010001100110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010001100110010) && ({row_reg, col_reg}<16'b0010001100110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010001100110100) && ({row_reg, col_reg}<16'b0010001100110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010001100110111) && ({row_reg, col_reg}<16'b0010001100111001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010001100111001) && ({row_reg, col_reg}<16'b0010001100111100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010001100111100) && ({row_reg, col_reg}<16'b0010001101000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001101000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001101000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001101000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010001101000111) && ({row_reg, col_reg}<16'b0010001101001001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010001101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001101001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001101001011) && ({row_reg, col_reg}<16'b0010001101001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010001101001101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010001101001110) && ({row_reg, col_reg}<16'b0010001101010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001101010000) && ({row_reg, col_reg}<16'b0010001101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010001101010101) && ({row_reg, col_reg}<16'b0010001101010111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010001101010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001101011000) && ({row_reg, col_reg}<16'b0010001101011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001101011111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010001101100000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010001101100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010001101100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001101100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001101100100)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b0010001101100101) && ({row_reg, col_reg}<16'b0010001101101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001101101000) && ({row_reg, col_reg}<16'b0010001101101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010001101101011) && ({row_reg, col_reg}<16'b0010001101101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001101101101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0010001101101110) && ({row_reg, col_reg}<16'b0010001101110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001101110000) && ({row_reg, col_reg}<16'b0010001101110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001101110010) && ({row_reg, col_reg}<16'b0010001101110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001101110111) && ({row_reg, col_reg}<16'b0010001101111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001101111001) && ({row_reg, col_reg}<16'b0010001101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010001101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001101111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010001101111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001101111110) && ({row_reg, col_reg}<16'b0010001110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001110000000) && ({row_reg, col_reg}<16'b0010001110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001110000011) && ({row_reg, col_reg}<16'b0010001110100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010001110100011) && ({row_reg, col_reg}<16'b0010001110101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001110101000) && ({row_reg, col_reg}<16'b0010001110101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001110101010) && ({row_reg, col_reg}<16'b0010001110101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001110101100) && ({row_reg, col_reg}<16'b0010001110101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010001110101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001110101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001110110000) && ({row_reg, col_reg}<16'b0010001110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010001110110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001110110100) && ({row_reg, col_reg}<16'b0010001110111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001110111010) && ({row_reg, col_reg}<16'b0010001111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001111000000) && ({row_reg, col_reg}<16'b0010001111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001111000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001111000110) && ({row_reg, col_reg}<16'b0010001111001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001111001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001111001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001111001011) && ({row_reg, col_reg}<16'b0010001111001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010001111001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001111001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001111001111) && ({row_reg, col_reg}<16'b0010001111010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010001111010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001111010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010001111010101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010001111010110) && ({row_reg, col_reg}<16'b0010001111011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001111011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010001111011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001111011101) && ({row_reg, col_reg}<16'b0010001111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001111011111) && ({row_reg, col_reg}<16'b0010001111100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001111100001) && ({row_reg, col_reg}<16'b0010001111100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001111100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001111100100) && ({row_reg, col_reg}<16'b0010001111101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001111101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001111101110) && ({row_reg, col_reg}<16'b0010001111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001111110010) && ({row_reg, col_reg}<16'b0010001111111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010001111111001) && ({row_reg, col_reg}<16'b0010001111111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0010001111111011) && ({row_reg, col_reg}<16'b0010010000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010000000000) && ({row_reg, col_reg}<16'b0010010000000011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010010000000011) && ({row_reg, col_reg}<16'b0010010000000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010000000101) && ({row_reg, col_reg}<16'b0010010000000111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010000000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010010000001000) && ({row_reg, col_reg}<16'b0010010000001010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010010000001010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010010000001011) && ({row_reg, col_reg}<16'b0010010000001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010000001111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010010000010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010000010010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010010000010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010010000010100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010010000010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010010000010110) && ({row_reg, col_reg}<16'b0010010000011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010000011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010000011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010010000011010) && ({row_reg, col_reg}<16'b0010010000011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010010000011100) && ({row_reg, col_reg}<16'b0010010000011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010010000011110) && ({row_reg, col_reg}<16'b0010010000100000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010010000100000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010010000100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010010000100010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0010010000100011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010010000100100)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0010010000100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010010000100110) && ({row_reg, col_reg}<16'b0010010000101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010010000101000) && ({row_reg, col_reg}<16'b0010010000101010)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0010010000101010) && ({row_reg, col_reg}<16'b0010010000101100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010000101100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010010000101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010000101110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010010000101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010010000110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010010000110001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0010010000110010) && ({row_reg, col_reg}<16'b0010010000110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010000110100) && ({row_reg, col_reg}<16'b0010010000111000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010000111000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010000111001)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010010000111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010000111011) && ({row_reg, col_reg}<16'b0010010000111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010000111101) && ({row_reg, col_reg}<16'b0010010001000001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010001000001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0010010001000010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010010001000011) && ({row_reg, col_reg}<16'b0010010001000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010001000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010001000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010001000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010010001001000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010010001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010010001001010) && ({row_reg, col_reg}<16'b0010010001001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010001001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010010001001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010001001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010001010000) && ({row_reg, col_reg}<16'b0010010001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010001010101) && ({row_reg, col_reg}<16'b0010010001010111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010010001010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010001011000) && ({row_reg, col_reg}<16'b0010010001011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010001011011) && ({row_reg, col_reg}<16'b0010010001011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010001011101) && ({row_reg, col_reg}<16'b0010010001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010001011111) && ({row_reg, col_reg}<16'b0010010001100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010010001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010001100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010010001100100)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b0010010001100101) && ({row_reg, col_reg}<16'b0010010001100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010001100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010010001101000) && ({row_reg, col_reg}<16'b0010010001101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010010001101010)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}>=16'b0010010001101011) && ({row_reg, col_reg}<16'b0010010001101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010001101101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0010010001101110) && ({row_reg, col_reg}<16'b0010010001110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010001110000) && ({row_reg, col_reg}<16'b0010010001110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010001110010) && ({row_reg, col_reg}<16'b0010010001111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010010001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010001111001) && ({row_reg, col_reg}<16'b0010010001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010010001111011) && ({row_reg, col_reg}<16'b0010010001111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010010001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010010000000) && ({row_reg, col_reg}<16'b0010010010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010010000011) && ({row_reg, col_reg}<16'b0010010010100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010010010100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010010100100) && ({row_reg, col_reg}<16'b0010010010101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010010101100) && ({row_reg, col_reg}<16'b0010010010101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010010101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010010010101111) && ({row_reg, col_reg}<16'b0010010010110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010010110001) && ({row_reg, col_reg}<16'b0010010010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010010010110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010010110100) && ({row_reg, col_reg}<16'b0010010010111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010010111010) && ({row_reg, col_reg}<16'b0010010011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010010011000000) && ({row_reg, col_reg}<16'b0010010011000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010011000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010011000110) && ({row_reg, col_reg}<16'b0010010011001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010011001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010011001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010011001011) && ({row_reg, col_reg}<16'b0010010011001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010010011001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010011001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010010011001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010011010000) && ({row_reg, col_reg}<16'b0010010011010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010010011010010) && ({row_reg, col_reg}<16'b0010010011010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010011010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010010011010101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010010011010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010011010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010010011011000) && ({row_reg, col_reg}<16'b0010010011011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010011011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010010011011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010010011011101) && ({row_reg, col_reg}<16'b0010010011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010011011111) && ({row_reg, col_reg}<16'b0010010011100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010011100001) && ({row_reg, col_reg}<16'b0010010011100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010011100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010011100100) && ({row_reg, col_reg}<16'b0010010011100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010011100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010011100111) && ({row_reg, col_reg}<16'b0010010011101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010011101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010010011101101) && ({row_reg, col_reg}<16'b0010010011110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010011110000) && ({row_reg, col_reg}<16'b0010010011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010011110010) && ({row_reg, col_reg}<16'b0010010011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010010011111001) && ({row_reg, col_reg}<16'b0010010011111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010011111011) && ({row_reg, col_reg}<16'b0010010011111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010011111101)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0010010011111110) && ({row_reg, col_reg}<16'b0010010100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010100000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010100000001) && ({row_reg, col_reg}<16'b0010010100000011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010010100000011) && ({row_reg, col_reg}<16'b0010010100000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010100000101) && ({row_reg, col_reg}<16'b0010010100000111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010100000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010010100001000) && ({row_reg, col_reg}<16'b0010010100001010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010010100001010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010010100001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010100001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010010100001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010010100001110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0010010100001111) && ({row_reg, col_reg}<16'b0010010100010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010100010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010010100010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010100010011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010010100010100) && ({row_reg, col_reg}<16'b0010010100010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010100010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010100010111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010010100011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010100011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010100011010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010010100011011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010010100011100) && ({row_reg, col_reg}<16'b0010010100011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010100011111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010010100100000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010010100100001) && ({row_reg, col_reg}<16'b0010010100100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010010100100101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0010010100100110) && ({row_reg, col_reg}<16'b0010010100101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010010100101000) && ({row_reg, col_reg}<16'b0010010100101010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010010100101010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010100101011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010010100101100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010100101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010010100101110) && ({row_reg, col_reg}<16'b0010010100110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010010100110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010010100110001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0010010100110010) && ({row_reg, col_reg}<16'b0010010100110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010100110100) && ({row_reg, col_reg}<16'b0010010100111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010010100111001) && ({row_reg, col_reg}<16'b0010010100111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010100111011) && ({row_reg, col_reg}<16'b0010010100111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010100111101) && ({row_reg, col_reg}<16'b0010010101000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010101000000) && ({row_reg, col_reg}<16'b0010010101000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010010101000011) && ({row_reg, col_reg}<16'b0010010101000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010101000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010101000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010010101000111) && ({row_reg, col_reg}<16'b0010010101001001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010010101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010010101001010) && ({row_reg, col_reg}<16'b0010010101001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010101001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010101001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010101001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010101010000) && ({row_reg, col_reg}<16'b0010010101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010101010101) && ({row_reg, col_reg}<16'b0010010101010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010101010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010010101011000) && ({row_reg, col_reg}<16'b0010010101011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010101011010) && ({row_reg, col_reg}<16'b0010010101011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010101011100) && ({row_reg, col_reg}<16'b0010010101011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010010101011110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010010101011111) && ({row_reg, col_reg}<16'b0010010101100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010010101100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010101100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010010101100100) && ({row_reg, col_reg}<16'b0010010101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010010101101100) && ({row_reg, col_reg}<16'b0010010101101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010010101101110) && ({row_reg, col_reg}<16'b0010010101110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010010101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010101110001) && ({row_reg, col_reg}<16'b0010010101111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010101111000) && ({row_reg, col_reg}<16'b0010010101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010101111011) && ({row_reg, col_reg}<16'b0010010101111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010010101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010110000000) && ({row_reg, col_reg}<16'b0010010110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010110000011) && ({row_reg, col_reg}<16'b0010010110100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010010110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010110100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010110100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010110100111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010110101000) && ({row_reg, col_reg}<16'b0010010110101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010110101100) && ({row_reg, col_reg}<16'b0010010110101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010110101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010110101111) && ({row_reg, col_reg}<16'b0010010110110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010010110110001) && ({row_reg, col_reg}<16'b0010010110110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010110110100) && ({row_reg, col_reg}<16'b0010010110111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010110111011) && ({row_reg, col_reg}<16'b0010010110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010010110111101) && ({row_reg, col_reg}<16'b0010010110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010010110111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010111000000) && ({row_reg, col_reg}<16'b0010010111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010111000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010111000110) && ({row_reg, col_reg}<16'b0010010111001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010111001011) && ({row_reg, col_reg}<16'b0010010111010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010111010010) && ({row_reg, col_reg}<16'b0010010111010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010111010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010010111010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010111010110) && ({row_reg, col_reg}<16'b0010010111011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010010111011000) && ({row_reg, col_reg}<16'b0010010111011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010111011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010010111011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010010111011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010111011101) && ({row_reg, col_reg}<16'b0010010111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010111011111) && ({row_reg, col_reg}<16'b0010010111100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010111100001) && ({row_reg, col_reg}<16'b0010010111100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010111100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010111100100) && ({row_reg, col_reg}<16'b0010010111101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010111101010) && ({row_reg, col_reg}<16'b0010010111101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010010111101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010111101110) && ({row_reg, col_reg}<16'b0010010111110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010111110000) && ({row_reg, col_reg}<16'b0010010111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010111110010) && ({row_reg, col_reg}<16'b0010010111111001)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0010010111111001) && ({row_reg, col_reg}<16'b0010011000000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010011000000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011000000001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010011000000010) && ({row_reg, col_reg}<16'b0010011000000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011000000101)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010011000000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010011000000111) && ({row_reg, col_reg}<16'b0010011000001011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010011000001011) && ({row_reg, col_reg}<16'b0010011000001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010011000001101) && ({row_reg, col_reg}<16'b0010011000010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010011000010001) && ({row_reg, col_reg}<16'b0010011000010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011000010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010011000010100) && ({row_reg, col_reg}<16'b0010011000010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010011000010110) && ({row_reg, col_reg}<16'b0010011000011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011000011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010011000011010) && ({row_reg, col_reg}<16'b0010011000011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010011000011100) && ({row_reg, col_reg}<16'b0010011000011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011000011111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0010011000100000) && ({row_reg, col_reg}<16'b0010011000100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010011000100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010011000100110) && ({row_reg, col_reg}<16'b0010011000101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011000101000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010011000101001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0010011000101010)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0010011000101011) && ({row_reg, col_reg}<16'b0010011000101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011000101101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0010011000101110) && ({row_reg, col_reg}<16'b0010011000110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010011000110000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010011000110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010011000110010) && ({row_reg, col_reg}<16'b0010011000110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010011000110100) && ({row_reg, col_reg}<16'b0010011000111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011000111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010011000111011) && ({row_reg, col_reg}<16'b0010011000111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011000111101) && ({row_reg, col_reg}<16'b0010011001000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010011001000000) && ({row_reg, col_reg}<16'b0010011001000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010011001000011) && ({row_reg, col_reg}<16'b0010011001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011001000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011001000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010011001000111) && ({row_reg, col_reg}<16'b0010011001001001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010011001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011001001011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0010011001001100) && ({row_reg, col_reg}<16'b0010011001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011001001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010011001010000) && ({row_reg, col_reg}<16'b0010011001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011001010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011001010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010011001010111)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0010011001011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011001011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011001011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011001011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010011001011100) && ({row_reg, col_reg}<16'b0010011001011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010011001011110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011001011111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010011001100000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010011001100001)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010011001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011001100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011001100100) && ({row_reg, col_reg}<16'b0010011001101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010011001101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010011001101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011001101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010011001101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010011001110000) && ({row_reg, col_reg}<16'b0010011001110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011001110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010011001110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010011001110100) && ({row_reg, col_reg}<16'b0010011001111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011001111000) && ({row_reg, col_reg}<16'b0010011001111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011001111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011001111011) && ({row_reg, col_reg}<16'b0010011001111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011010000000) && ({row_reg, col_reg}<16'b0010011010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011010000011) && ({row_reg, col_reg}<16'b0010011010100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010011010100100) && ({row_reg, col_reg}<16'b0010011010100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010011010100111) && ({row_reg, col_reg}<16'b0010011010101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011010101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010011010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011010101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011010101111) && ({row_reg, col_reg}<16'b0010011010110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010011010110001) && ({row_reg, col_reg}<16'b0010011010110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011010110100) && ({row_reg, col_reg}<16'b0010011010111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011010111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010011010111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011010111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010011010111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010011011000000) && ({row_reg, col_reg}<16'b0010011011000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011011000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010011011000110) && ({row_reg, col_reg}<16'b0010011011001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011011001011) && ({row_reg, col_reg}<16'b0010011011001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010011011001101) && ({row_reg, col_reg}<16'b0010011011010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011011010000) && ({row_reg, col_reg}<16'b0010011011010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011011010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011011010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010011011010101) && ({row_reg, col_reg}<16'b0010011011011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011011011010) && ({row_reg, col_reg}<16'b0010011011011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010011011011100) && ({row_reg, col_reg}<16'b0010011011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011011011111) && ({row_reg, col_reg}<16'b0010011011100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010011011100001) && ({row_reg, col_reg}<16'b0010011011100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011011100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011011100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010011011100101) && ({row_reg, col_reg}<16'b0010011011101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011011101001) && ({row_reg, col_reg}<16'b0010011011101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010011011101011) && ({row_reg, col_reg}<16'b0010011011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011011110010) && ({row_reg, col_reg}<16'b0010011011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011011111001)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0010011011111010) && ({row_reg, col_reg}<16'b0010011100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010011100000000) && ({row_reg, col_reg}<16'b0010011100000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010011100000010) && ({row_reg, col_reg}<16'b0010011100000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011100000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011100000111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010011100001000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0010011100001001) && ({row_reg, col_reg}<16'b0010011100001011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010011100001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011100001100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011100001101)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010011100001110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010011100001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011100010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010011100010001) && ({row_reg, col_reg}<16'b0010011100010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010011100010011) && ({row_reg, col_reg}<16'b0010011100010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010011100010101) && ({row_reg, col_reg}<16'b0010011100011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011100011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011100011001)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0010011100011010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010011100011011) && ({row_reg, col_reg}<16'b0010011100011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011100011101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010011100011110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010011100011111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0010011100100000) && ({row_reg, col_reg}<16'b0010011100100010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010011100100010)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0010011100100011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010011100100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010011100100101) && ({row_reg, col_reg}<16'b0010011100100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011100100111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010011100101000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010011100101001) && ({row_reg, col_reg}<16'b0010011100101011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0010011100101011) && ({row_reg, col_reg}<16'b0010011100101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011100101101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0010011100101110) && ({row_reg, col_reg}<16'b0010011100110001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010011100110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011100110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011100110011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010011100110100) && ({row_reg, col_reg}<16'b0010011100110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011100110110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010011100110111) && ({row_reg, col_reg}<16'b0010011100111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011100111010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010011100111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011100111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011100111101) && ({row_reg, col_reg}<16'b0010011101000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010011101000000) && ({row_reg, col_reg}<16'b0010011101000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010011101000011) && ({row_reg, col_reg}<16'b0010011101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010011101000101) && ({row_reg, col_reg}<16'b0010011101001010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010011101001011) && ({row_reg, col_reg}<16'b0010011101001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011101001110) && ({row_reg, col_reg}<16'b0010011101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010011101010000) && ({row_reg, col_reg}<16'b0010011101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010011101010100) && ({row_reg, col_reg}<16'b0010011101010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011101010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011101010111) && ({row_reg, col_reg}<16'b0010011101011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011101011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010011101011010) && ({row_reg, col_reg}<16'b0010011101011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011101011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011101011110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0010011101011111) && ({row_reg, col_reg}<16'b0010011101100010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011101100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010011101100100) && ({row_reg, col_reg}<16'b0010011101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010011101101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010011101101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011101101110) && ({row_reg, col_reg}<16'b0010011101110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010011101110000) && ({row_reg, col_reg}<16'b0010011101110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010011101110010) && ({row_reg, col_reg}<16'b0010011101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010011101110100) && ({row_reg, col_reg}<16'b0010011101111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011101111000) && ({row_reg, col_reg}<16'b0010011101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011101111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011101111100) && ({row_reg, col_reg}<16'b0010011101111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011110000000) && ({row_reg, col_reg}<16'b0010011110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011110000011) && ({row_reg, col_reg}<16'b0010011110100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011110100101) && ({row_reg, col_reg}<16'b0010011110100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010011110100111) && ({row_reg, col_reg}<16'b0010011110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011110101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010011110101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011110101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011110101101) && ({row_reg, col_reg}<16'b0010011110101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010011110101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011110110000) && ({row_reg, col_reg}<16'b0010011110110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010011110110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010011110110110) && ({row_reg, col_reg}<16'b0010011110111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011110111010) && ({row_reg, col_reg}<16'b0010011110111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011110111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010011110111101) && ({row_reg, col_reg}<16'b0010011110111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011110111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010011111000000) && ({row_reg, col_reg}<16'b0010011111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011111000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010011111000110) && ({row_reg, col_reg}<16'b0010011111001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011111001011) && ({row_reg, col_reg}<16'b0010011111001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011111001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011111001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010011111001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011111010000) && ({row_reg, col_reg}<16'b0010011111010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010011111010010) && ({row_reg, col_reg}<16'b0010011111010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011111010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010011111010101) && ({row_reg, col_reg}<16'b0010011111011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011111011010) && ({row_reg, col_reg}<16'b0010011111011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011111011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011111011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010011111011110) && ({row_reg, col_reg}<16'b0010011111100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011111100010) && ({row_reg, col_reg}<16'b0010011111101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010011111101001) && ({row_reg, col_reg}<16'b0010011111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011111101111) && ({row_reg, col_reg}<16'b0010011111110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010011111110001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0010011111110010) && ({row_reg, col_reg}<16'b0010100000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100000000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100000000001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010100000000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100000000011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0010100000000100) && ({row_reg, col_reg}<16'b0010100000000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100000000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100000000111) && ({row_reg, col_reg}<16'b0010100000001011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010100000001011) && ({row_reg, col_reg}<16'b0010100000010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100000010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010100000010001) && ({row_reg, col_reg}<16'b0010100000010011)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}>=16'b0010100000010011) && ({row_reg, col_reg}<16'b0010100000010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010100000010101) && ({row_reg, col_reg}<16'b0010100000011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100000011001)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0010100000011010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010100000011011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010100000011100) && ({row_reg, col_reg}<16'b0010100000011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100000011110)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0010100000011111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0010100000100000) && ({row_reg, col_reg}<16'b0010100000100010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010100000100010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0010100000100011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010100000100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010100000100101) && ({row_reg, col_reg}<16'b0010100000101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100000101000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010100000101001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0010100000101010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0010100000101011) && ({row_reg, col_reg}<16'b0010100000101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010100000101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100000101110) && ({row_reg, col_reg}<16'b0010100000110001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010100000110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100000110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100000110011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010100000110100) && ({row_reg, col_reg}<16'b0010100000110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100000110110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010100000110111) && ({row_reg, col_reg}<16'b0010100000111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100000111011) && ({row_reg, col_reg}<16'b0010100000111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100000111101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010100000111110) && ({row_reg, col_reg}<16'b0010100001000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100001000001) && ({row_reg, col_reg}<16'b0010100001000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010100001000011) && ({row_reg, col_reg}<16'b0010100001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010100001000101) && ({row_reg, col_reg}<16'b0010100001001010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100001001010) && ({row_reg, col_reg}<16'b0010100001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010100001010000) && ({row_reg, col_reg}<16'b0010100001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010100001010100) && ({row_reg, col_reg}<16'b0010100001011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010100001011000) && ({row_reg, col_reg}<16'b0010100001011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010100001011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100001011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010100001011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010100001011101) && ({row_reg, col_reg}<16'b0010100001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010100001011111) && ({row_reg, col_reg}<16'b0010100001100010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010100001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100001100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010100001100100) && ({row_reg, col_reg}<16'b0010100001101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100001101100) && ({row_reg, col_reg}<16'b0010100001110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010100001110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010100001110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100001110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010100001110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100001110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010100001110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010100001110110) && ({row_reg, col_reg}<16'b0010100001111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100001111000) && ({row_reg, col_reg}<16'b0010100001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100001111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010100001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100001111110) && ({row_reg, col_reg}<16'b0010100010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100010000000) && ({row_reg, col_reg}<16'b0010100010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100010000011) && ({row_reg, col_reg}<16'b0010100010100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100010100101) && ({row_reg, col_reg}<16'b0010100010100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100010100111) && ({row_reg, col_reg}<16'b0010100010101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100010101011) && ({row_reg, col_reg}<16'b0010100010101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100010101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100010110000) && ({row_reg, col_reg}<16'b0010100010110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100010110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010100010110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100010110100) && ({row_reg, col_reg}<16'b0010100010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100010110110) && ({row_reg, col_reg}<16'b0010100010111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100010111010) && ({row_reg, col_reg}<16'b0010100010111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010100010111100) && ({row_reg, col_reg}<16'b0010100010111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100010111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010100011000000) && ({row_reg, col_reg}<16'b0010100011000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100011000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100011000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010100011000111) && ({row_reg, col_reg}<16'b0010100011001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100011001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010100011001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100011001101) && ({row_reg, col_reg}<16'b0010100011001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010100011001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100011010000) && ({row_reg, col_reg}<16'b0010100011010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010100011010010) && ({row_reg, col_reg}<16'b0010100011010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100011010100) && ({row_reg, col_reg}<16'b0010100011010110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010100011010110) && ({row_reg, col_reg}<16'b0010100011011000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0010100011011000) && ({row_reg, col_reg}<16'b0010100011011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100011011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010100011011011) && ({row_reg, col_reg}<16'b0010100011011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100011011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100011011110) && ({row_reg, col_reg}<16'b0010100011101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100011101010) && ({row_reg, col_reg}<16'b0010100011101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010100011101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100011101111) && ({row_reg, col_reg}<16'b0010100011110010)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0010100011110010) && ({row_reg, col_reg}<16'b0010100100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100100000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010100100000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100100000010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0010100100000011) && ({row_reg, col_reg}<16'b0010100100000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010100100000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100100000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100100000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010100100001000) && ({row_reg, col_reg}<16'b0010100100001010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010100100001010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010100100001011) && ({row_reg, col_reg}<16'b0010100100001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100100001110) && ({row_reg, col_reg}<16'b0010100100010000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010100100010000) && ({row_reg, col_reg}<16'b0010100100010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010100100010010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010100100010011) && ({row_reg, col_reg}<16'b0010100100010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010100100010101) && ({row_reg, col_reg}<16'b0010100100011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100100011010) && ({row_reg, col_reg}<16'b0010100100011100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010100100011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010100100011101) && ({row_reg, col_reg}<16'b0010100100100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100100100000) && ({row_reg, col_reg}<16'b0010100100100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010100100100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100100100110) && ({row_reg, col_reg}<16'b0010100100101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010100100101000) && ({row_reg, col_reg}<16'b0010100100101010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010100100101010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100100101011) && ({row_reg, col_reg}<16'b0010100100101110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010100100101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100100101111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010100100110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010100100110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100100110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100100110011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010100100110100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100100110101) && ({row_reg, col_reg}<16'b0010100100110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010100100110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100100111000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010100100111001) && ({row_reg, col_reg}<16'b0010100100111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100100111011) && ({row_reg, col_reg}<16'b0010100100111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100100111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100100111110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010100100111111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010100101000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100101000001) && ({row_reg, col_reg}<16'b0010100101000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010100101000011) && ({row_reg, col_reg}<16'b0010100101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100101000101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010100101000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100101000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010100101001000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010100101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100101001010) && ({row_reg, col_reg}<16'b0010100101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010100101001100) && ({row_reg, col_reg}<16'b0010100101001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100101001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010100101001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100101010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010100101010001) && ({row_reg, col_reg}<16'b0010100101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010100101010100) && ({row_reg, col_reg}<16'b0010100101010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010100101010111) && ({row_reg, col_reg}<16'b0010100101011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010100101011101) && ({row_reg, col_reg}<16'b0010100101100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100101100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010100101100100) && ({row_reg, col_reg}<16'b0010100101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100101101100) && ({row_reg, col_reg}<16'b0010100101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100101101110) && ({row_reg, col_reg}<16'b0010100101110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100101110000) && ({row_reg, col_reg}<16'b0010100101110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100101110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010100101110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100101110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010100101110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100101110111) && ({row_reg, col_reg}<16'b0010100101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100110000000) && ({row_reg, col_reg}<16'b0010100110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100110000011) && ({row_reg, col_reg}<16'b0010100110100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010100110100100) && ({row_reg, col_reg}<16'b0010100110100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100110100110) && ({row_reg, col_reg}<16'b0010100110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100110101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100110101100) && ({row_reg, col_reg}<16'b0010100110101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010100110101110) && ({row_reg, col_reg}<16'b0010100110110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100110110000) && ({row_reg, col_reg}<16'b0010100110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010100110110011) && ({row_reg, col_reg}<16'b0010100110110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100110110110) && ({row_reg, col_reg}<16'b0010100110111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100110111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010100110111011) && ({row_reg, col_reg}<16'b0010100111000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010100111000000) && ({row_reg, col_reg}<16'b0010100111000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100111000110) && ({row_reg, col_reg}<16'b0010100111001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010100111001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100111001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010100111001011) && ({row_reg, col_reg}<16'b0010100111001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010100111001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100111010000) && ({row_reg, col_reg}<16'b0010100111010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010100111010010) && ({row_reg, col_reg}<16'b0010100111010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100111010101) && ({row_reg, col_reg}<16'b0010100111011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010100111011010) && ({row_reg, col_reg}<16'b0010100111011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100111011101) && ({row_reg, col_reg}<16'b0010100111100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100111100001) && ({row_reg, col_reg}<16'b0010100111100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100111100101) && ({row_reg, col_reg}<16'b0010100111101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100111101100) && ({row_reg, col_reg}<16'b0010100111110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100111110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010100111110001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0010100111110010) && ({row_reg, col_reg}<16'b0010101000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010101000000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010101000000001) && ({row_reg, col_reg}<16'b0010101000000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101000000011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0010101000000100) && ({row_reg, col_reg}<16'b0010101000000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101000000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101000000111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010101000001000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101000001001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0010101000001010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010101000001011) && ({row_reg, col_reg}<16'b0010101000001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010101000001110) && ({row_reg, col_reg}<16'b0010101000010000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010101000010000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010101000010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101000010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010101000010011) && ({row_reg, col_reg}<16'b0010101000010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010101000010101) && ({row_reg, col_reg}<16'b0010101000011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010101000011011) && ({row_reg, col_reg}<16'b0010101000011101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010101000011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101000011110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010101000011111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010101000100000) && ({row_reg, col_reg}<16'b0010101000100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101000100100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010101000100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010101000100110) && ({row_reg, col_reg}<16'b0010101000101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010101000101000) && ({row_reg, col_reg}<16'b0010101000101010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010101000101010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010101000101011) && ({row_reg, col_reg}<16'b0010101000101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101000101101)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010101000101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101000101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010101000110000) && ({row_reg, col_reg}<16'b0010101000110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010101000110010) && ({row_reg, col_reg}<16'b0010101000110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101000110100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010101000110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101000110110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010101000110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101000111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101000111001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010101000111010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0010101000111011) && ({row_reg, col_reg}<16'b0010101000111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101000111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101000111110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010101000111111) && ({row_reg, col_reg}<16'b0010101001000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010101001000001) && ({row_reg, col_reg}<16'b0010101001000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010101001000011) && ({row_reg, col_reg}<16'b0010101001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101001000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010101001000111) && ({row_reg, col_reg}<16'b0010101001001001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010101001001010) && ({row_reg, col_reg}<16'b0010101001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101001001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010101001001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101001001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010101001001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101001010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010101001010001) && ({row_reg, col_reg}<16'b0010101001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010101001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010101001010101) && ({row_reg, col_reg}<16'b0010101001011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010101001011000) && ({row_reg, col_reg}<16'b0010101001011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101001011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010101001011100) && ({row_reg, col_reg}<16'b0010101001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101001100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010101001100011) && ({row_reg, col_reg}<16'b0010101001101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101001101100) && ({row_reg, col_reg}<16'b0010101001110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101001110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010101001110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010101001110100) && ({row_reg, col_reg}<16'b0010101001110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101001110111) && ({row_reg, col_reg}<16'b0010101001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101010000000) && ({row_reg, col_reg}<16'b0010101010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101010000011) && ({row_reg, col_reg}<16'b0010101010100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010101010100100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101010100101) && ({row_reg, col_reg}<16'b0010101010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101010101101) && ({row_reg, col_reg}<16'b0010101010101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101010101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101010110000) && ({row_reg, col_reg}<16'b0010101010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010101010110011) && ({row_reg, col_reg}<16'b0010101010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101010110101) && ({row_reg, col_reg}<16'b0010101010111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101010111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010101010111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101010111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010101010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101010111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010101011000000) && ({row_reg, col_reg}<16'b0010101011000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101011000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010101011000110) && ({row_reg, col_reg}<16'b0010101011001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010101011001000) && ({row_reg, col_reg}<16'b0010101011001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101011001100) && ({row_reg, col_reg}<16'b0010101011010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101011010000) && ({row_reg, col_reg}<16'b0010101011010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010101011010010) && ({row_reg, col_reg}<16'b0010101011011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101011011101) && ({row_reg, col_reg}<16'b0010101011100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101011100010) && ({row_reg, col_reg}<16'b0010101011100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101011100100) && ({row_reg, col_reg}<16'b0010101011100110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101011100110) && ({row_reg, col_reg}<16'b0010101011101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010101011101000) && ({row_reg, col_reg}<16'b0010101011101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101011101100) && ({row_reg, col_reg}<16'b0010101011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101011101111) && ({row_reg, col_reg}<16'b0010101011110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101011110001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0010101011110010) && ({row_reg, col_reg}<16'b0010101100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010101100000000) && ({row_reg, col_reg}<16'b0010101100000010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010101100000010) && ({row_reg, col_reg}<16'b0010101100000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101100000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101100000111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010101100001000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0010101100001001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010101100001010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101100001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010101100001100) && ({row_reg, col_reg}<16'b0010101100001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010101100001110) && ({row_reg, col_reg}<16'b0010101100010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101100010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101100010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101100010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010101100010011) && ({row_reg, col_reg}<16'b0010101100010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010101100010101) && ({row_reg, col_reg}<16'b0010101100010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010101100010111) && ({row_reg, col_reg}<16'b0010101100011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010101100011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101100011011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010101100011100) && ({row_reg, col_reg}<16'b0010101100011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101100011110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010101100011111) && ({row_reg, col_reg}<16'b0010101100100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101100100001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010101100100010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010101100100011) && ({row_reg, col_reg}<16'b0010101100100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010101100100101) && ({row_reg, col_reg}<16'b0010101100100111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010101100100111) && ({row_reg, col_reg}<16'b0010101100101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101100101001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010101100101010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0010101100101011) && ({row_reg, col_reg}<16'b0010101100101110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010101100101110) && ({row_reg, col_reg}<16'b0010101100110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101100110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010101100110011) && ({row_reg, col_reg}<16'b0010101100110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101100110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101100111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101100111001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010101100111010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010101100111011) && ({row_reg, col_reg}<16'b0010101100111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010101100111101) && ({row_reg, col_reg}<16'b0010101100111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101100111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010101101000000) && ({row_reg, col_reg}<16'b0010101101000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010101101000011) && ({row_reg, col_reg}<16'b0010101101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101101000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010101101000111) && ({row_reg, col_reg}<16'b0010101101001001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010101101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010101101001010) && ({row_reg, col_reg}<16'b0010101101001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101101001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010101101001110) && ({row_reg, col_reg}<16'b0010101101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101101010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010101101010001) && ({row_reg, col_reg}<16'b0010101101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010101101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010101101010101) && ({row_reg, col_reg}<16'b0010101101010111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010101101010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010101101011000) && ({row_reg, col_reg}<16'b0010101101100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010101101100011) && ({row_reg, col_reg}<16'b0010101101100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101101100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010101101100110) && ({row_reg, col_reg}<16'b0010101101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101101101100) && ({row_reg, col_reg}<16'b0010101101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101101101110) && ({row_reg, col_reg}<16'b0010101101110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010101101110000) && ({row_reg, col_reg}<16'b0010101101110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101101110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010101101110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010101101110100) && ({row_reg, col_reg}<16'b0010101101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101101110110) && ({row_reg, col_reg}<16'b0010101101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101101111011) && ({row_reg, col_reg}<16'b0010101101111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101101111101) && ({row_reg, col_reg}<16'b0010101101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101110000000) && ({row_reg, col_reg}<16'b0010101110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101110000011) && ({row_reg, col_reg}<16'b0010101110100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010101110100100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101110100101) && ({row_reg, col_reg}<16'b0010101110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101110101001) && ({row_reg, col_reg}<16'b0010101110101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101110101011) && ({row_reg, col_reg}<16'b0010101110101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101110101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101110110000) && ({row_reg, col_reg}<16'b0010101110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010101110110011) && ({row_reg, col_reg}<16'b0010101110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101110110101) && ({row_reg, col_reg}<16'b0010101110111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101110111001) && ({row_reg, col_reg}<16'b0010101110111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101110111100) && ({row_reg, col_reg}<16'b0010101111000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010101111000000) && ({row_reg, col_reg}<16'b0010101111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101111000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010101111000110) && ({row_reg, col_reg}<16'b0010101111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101111001011) && ({row_reg, col_reg}<16'b0010101111010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101111010000) && ({row_reg, col_reg}<16'b0010101111010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010101111010011) && ({row_reg, col_reg}<16'b0010101111011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101111011000) && ({row_reg, col_reg}<16'b0010101111011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010101111011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010101111011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101111011100) && ({row_reg, col_reg}<16'b0010101111100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101111100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101111100001) && ({row_reg, col_reg}<16'b0010101111100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101111100011) && ({row_reg, col_reg}<16'b0010101111100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101111100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010101111100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010101111100111) && ({row_reg, col_reg}<16'b0010101111101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101111101001) && ({row_reg, col_reg}<16'b0010101111101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101111101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101111101100) && ({row_reg, col_reg}<16'b0010101111101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101111101110) && ({row_reg, col_reg}<16'b0010101111110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101111110001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0010101111110010) && ({row_reg, col_reg}<16'b0010110000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010110000000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010110000000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110000000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010110000000011) && ({row_reg, col_reg}<16'b0010110000000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110000000110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010110000000111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010110000001000) && ({row_reg, col_reg}<16'b0010110000001010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010110000001010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010110000001011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010110000001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110000001101)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=16'b0010110000001110) && ({row_reg, col_reg}<16'b0010110000010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010110000010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010110000010001) && ({row_reg, col_reg}<16'b0010110000010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010110000010011) && ({row_reg, col_reg}<16'b0010110000010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010110000010101) && ({row_reg, col_reg}<16'b0010110000010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010110000010111) && ({row_reg, col_reg}<16'b0010110000011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110000011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110000011010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010110000011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110000011100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==16'b0010110000011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110000011110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010110000011111) && ({row_reg, col_reg}<16'b0010110000100001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010110000100001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010110000100010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010110000100011) && ({row_reg, col_reg}<16'b0010110000100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010110000100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010110000100110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010110000100111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010110000101000)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0010110000101001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010110000101010) && ({row_reg, col_reg}<16'b0010110000101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110000101100)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}==16'b0010110000101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110000101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010110000101111) && ({row_reg, col_reg}<16'b0010110000110001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010110000110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110000110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010110000110011) && ({row_reg, col_reg}<16'b0010110000110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110000110101)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}==16'b0010110000110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110000110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110000111000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010110000111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110000111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010110000111011) && ({row_reg, col_reg}<16'b0010110000111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010110000111101) && ({row_reg, col_reg}<16'b0010110000111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110000111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010110001000000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0010110001000001) && ({row_reg, col_reg}<16'b0010110001000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010110001000011) && ({row_reg, col_reg}<16'b0010110001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110001000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010110001000111) && ({row_reg, col_reg}<16'b0010110001001001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010110001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010110001001100) && ({row_reg, col_reg}<16'b0010110001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010110001010000) && ({row_reg, col_reg}<16'b0010110001010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010110001010010)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0010110001010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010110001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110001010101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010110001010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110001010111) && ({row_reg, col_reg}<16'b0010110001011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010110001011001) && ({row_reg, col_reg}<16'b0010110001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110001100010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010110001100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110001100100)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==16'b0010110001100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010110001100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010110001100111) && ({row_reg, col_reg}<16'b0010110001101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110001101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110001101110) && ({row_reg, col_reg}<16'b0010110001110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010110001110000) && ({row_reg, col_reg}<16'b0010110001110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110001110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010110001110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110001110100) && ({row_reg, col_reg}<16'b0010110001110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110001110110) && ({row_reg, col_reg}<16'b0010110001111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110001111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110001111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110001111100) && ({row_reg, col_reg}<16'b0010110010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110010000000) && ({row_reg, col_reg}<16'b0010110010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110010000011) && ({row_reg, col_reg}<16'b0010110010100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010110010100100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110010100101) && ({row_reg, col_reg}<16'b0010110010100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110010100111) && ({row_reg, col_reg}<16'b0010110010101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010110010101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110010101011) && ({row_reg, col_reg}<16'b0010110010101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110010101110) && ({row_reg, col_reg}<16'b0010110010110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110010110000) && ({row_reg, col_reg}<16'b0010110010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110010110011) && ({row_reg, col_reg}<16'b0010110010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110010110101) && ({row_reg, col_reg}<16'b0010110011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110011001000) && ({row_reg, col_reg}<16'b0010110011001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010110011001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110011001011) && ({row_reg, col_reg}<16'b0010110011001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110011001101) && ({row_reg, col_reg}<16'b0010110011010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010110011010001) && ({row_reg, col_reg}<16'b0010110011010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110011010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010110011010100) && ({row_reg, col_reg}<16'b0010110011010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110011010110) && ({row_reg, col_reg}<16'b0010110011011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110011011100) && ({row_reg, col_reg}<16'b0010110011100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110011100100) && ({row_reg, col_reg}<16'b0010110011101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110011101110) && ({row_reg, col_reg}<16'b0010110011110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110011110001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0010110011110010) && ({row_reg, col_reg}<16'b0010110100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010110100000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010110100000001) && ({row_reg, col_reg}<16'b0010110100000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010110100000011) && ({row_reg, col_reg}<16'b0010110100000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110100000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110100000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010110100001000) && ({row_reg, col_reg}<16'b0010110100001010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010110100001010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0010110100001011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010110100001100) && ({row_reg, col_reg}<16'b0010110100010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110100010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010110100010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010110100010010) && ({row_reg, col_reg}<16'b0010110100010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010110100010101) && ({row_reg, col_reg}<16'b0010110100010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110100010111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010110100011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110100011001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010110100011010) && ({row_reg, col_reg}<16'b0010110100011111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010110100011111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010110100100000) && ({row_reg, col_reg}<16'b0010110100100010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010110100100010) && ({row_reg, col_reg}<16'b0010110100100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010110100100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010110100100110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010110100100111)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}>=16'b0010110100101000) && ({row_reg, col_reg}<16'b0010110100101010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0010110100101010)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0010110100101011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110100101100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010110100101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110100101110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010110100101111) && ({row_reg, col_reg}<16'b0010110100110001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010110100110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110100110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010110100110011) && ({row_reg, col_reg}<16'b0010110100110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110100110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110100110111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010110100111000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0010110100111001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010110100111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110100111011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010110100111100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110100111101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010110100111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110100111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010110101000000) && ({row_reg, col_reg}<16'b0010110101000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010110101000011) && ({row_reg, col_reg}<16'b0010110101000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110101000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010110101000111) && ({row_reg, col_reg}<16'b0010110101001001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010110101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110101001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010110101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010110101001100) && ({row_reg, col_reg}<16'b0010110101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010110101010000) && ({row_reg, col_reg}<16'b0010110101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010110101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010110101010101) && ({row_reg, col_reg}<16'b0010110101010111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110101010111) && ({row_reg, col_reg}<16'b0010110101011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010110101011001) && ({row_reg, col_reg}<16'b0010110101011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110101011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010110101100000) && ({row_reg, col_reg}<16'b0010110101100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110101100010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110101100011) && ({row_reg, col_reg}<16'b0010110101100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110101100101) && ({row_reg, col_reg}<16'b0010110101101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010110101101000) && ({row_reg, col_reg}<16'b0010110101101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110101101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110101101110) && ({row_reg, col_reg}<16'b0010110101110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010110101110000) && ({row_reg, col_reg}<16'b0010110101110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110101110010) && ({row_reg, col_reg}<16'b0010110101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110101110100) && ({row_reg, col_reg}<16'b0010110101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110101110110) && ({row_reg, col_reg}<16'b0010110101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110101111000) && ({row_reg, col_reg}<16'b0010110101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110101111011) && ({row_reg, col_reg}<16'b0010110110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110110000000) && ({row_reg, col_reg}<16'b0010110110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110110000011) && ({row_reg, col_reg}<16'b0010110110100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110110100100) && ({row_reg, col_reg}<16'b0010110110100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110110100111) && ({row_reg, col_reg}<16'b0010110110101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110110101010) && ({row_reg, col_reg}<16'b0010110110101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010110110101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010110110101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010110110101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110110110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110110110001) && ({row_reg, col_reg}<16'b0010110110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010110110110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110110110100) && ({row_reg, col_reg}<16'b0010110110110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110110110110) && ({row_reg, col_reg}<16'b0010110111000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110111000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110111000101) && ({row_reg, col_reg}<16'b0010110111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110111000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110111001000) && ({row_reg, col_reg}<16'b0010110111001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110111001010) && ({row_reg, col_reg}<16'b0010110111001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110111001100) && ({row_reg, col_reg}<16'b0010110111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110111001110) && ({row_reg, col_reg}<16'b0010110111010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010110111010001) && ({row_reg, col_reg}<16'b0010110111010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110111010110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110111010111) && ({row_reg, col_reg}<16'b0010110111011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110111011101) && ({row_reg, col_reg}<16'b0010110111100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110111100011) && ({row_reg, col_reg}<16'b0010110111101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110111101110) && ({row_reg, col_reg}<16'b0010110111110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110111110001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0010110111110010) && ({row_reg, col_reg}<16'b0010111000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010111000000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010111000000001) && ({row_reg, col_reg}<16'b0010111000000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010111000000100) && ({row_reg, col_reg}<16'b0010111000000110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010111000000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111000000111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0010111000001000) && ({row_reg, col_reg}<16'b0010111000001010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010111000001010)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0010111000001011)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=16'b0010111000001100) && ({row_reg, col_reg}<16'b0010111000001110)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0010111000001110)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0010111000001111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010111000010000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010111000010001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010111000010010) && ({row_reg, col_reg}<16'b0010111000010100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010111000010100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0010111000010101) && ({row_reg, col_reg}<16'b0010111000010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111000010111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010111000011000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010111000011001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010111000011010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0010111000011011)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0010111000011100)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==16'b0010111000011101)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==16'b0010111000011110)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0010111000011111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010111000100000) && ({row_reg, col_reg}<16'b0010111000100010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0010111000100010) && ({row_reg, col_reg}<16'b0010111000100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010111000100100) && ({row_reg, col_reg}<16'b0010111000100111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010111000100111)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0010111000101000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0010111000101001)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0010111000101010)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==16'b0010111000101011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0010111000101100) && ({row_reg, col_reg}<16'b0010111000101110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010111000101110) && ({row_reg, col_reg}<16'b0010111000110000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0010111000110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010111000110001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0010111000110010) && ({row_reg, col_reg}<16'b0010111000110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111000110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010111000110110)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0010111000110111)) color_data = 12'b100110000110;
		if(({row_reg, col_reg}==16'b0010111000111000)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0010111000111001)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0010111000111010)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0010111000111011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0010111000111100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0010111000111101) && ({row_reg, col_reg}<16'b0010111001000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010111001000011) && ({row_reg, col_reg}<16'b0010111001000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111001000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010111001000111) && ({row_reg, col_reg}<16'b0010111001001001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010111001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111001001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010111001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111001001100) && ({row_reg, col_reg}<16'b0010111001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010111001010000) && ({row_reg, col_reg}<16'b0010111001010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010111001010011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0010111001010100) && ({row_reg, col_reg}<16'b0010111001010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010111001010110) && ({row_reg, col_reg}<16'b0010111001011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111001011001) && ({row_reg, col_reg}<16'b0010111001011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010111001011110) && ({row_reg, col_reg}<16'b0010111001100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111001100000) && ({row_reg, col_reg}<16'b0010111001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111001100010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010111001100011) && ({row_reg, col_reg}<16'b0010111001100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111001100101) && ({row_reg, col_reg}<16'b0010111001101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010111001101000) && ({row_reg, col_reg}<16'b0010111001101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111001101100) && ({row_reg, col_reg}<16'b0010111001101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010111001101110) && ({row_reg, col_reg}<16'b0010111001110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111001110000) && ({row_reg, col_reg}<16'b0010111001110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111001110010) && ({row_reg, col_reg}<16'b0010111001110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010111001110100) && ({row_reg, col_reg}<16'b0010111001110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111001110110) && ({row_reg, col_reg}<16'b0010111001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111001111000) && ({row_reg, col_reg}<16'b0010111001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111001111100) && ({row_reg, col_reg}<16'b0010111010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111010000000) && ({row_reg, col_reg}<16'b0010111010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111010000011) && ({row_reg, col_reg}<16'b0010111010100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010111010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111010100101) && ({row_reg, col_reg}<16'b0010111010101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111010101000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=16'b0010111010101001) && ({row_reg, col_reg}<16'b0010111010101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010111010101011) && ({row_reg, col_reg}<16'b0010111010101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010111010101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010111010101110) && ({row_reg, col_reg}<16'b0010111010110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111010110001) && ({row_reg, col_reg}<16'b0010111010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010111010110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111010110100) && ({row_reg, col_reg}<16'b0010111010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111010110111) && ({row_reg, col_reg}<16'b0010111010111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111010111010) && ({row_reg, col_reg}<16'b0010111010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111010111110) && ({row_reg, col_reg}<16'b0010111011000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111011000000) && ({row_reg, col_reg}<16'b0010111011000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111011000011) && ({row_reg, col_reg}<16'b0010111011000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111011000101) && ({row_reg, col_reg}<16'b0010111011000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111011000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111011001000) && ({row_reg, col_reg}<16'b0010111011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010111011001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111011001100) && ({row_reg, col_reg}<16'b0010111011001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111011001111) && ({row_reg, col_reg}<16'b0010111011010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111011010001) && ({row_reg, col_reg}<16'b0010111011011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111011011110) && ({row_reg, col_reg}<16'b0010111011100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111011100010) && ({row_reg, col_reg}<16'b0010111011100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111011100100) && ({row_reg, col_reg}<16'b0010111011100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111011100110) && ({row_reg, col_reg}<16'b0010111011101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111011101011) && ({row_reg, col_reg}<16'b0010111011101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010111011101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111011101110) && ({row_reg, col_reg}<16'b0010111011110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111011110001)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0010111011110010) && ({row_reg, col_reg}<16'b0010111100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010111100000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111100000001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010111100000010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010111100000011) && ({row_reg, col_reg}<16'b0010111100000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010111100000101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0010111100000110) && ({row_reg, col_reg}<16'b0010111100001000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010111100001000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0010111100001001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010111100001010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0010111100001011)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0010111100001100)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0010111100001101)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==16'b0010111100001110)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0010111100001111)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0010111100010000)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}>=16'b0010111100010001) && ({row_reg, col_reg}<16'b0010111100010100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010111100010100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0010111100010101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010111100010110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010111100010111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010111100011000)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0010111100011001)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0010111100011010)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0010111100011011)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0010111100011100)) color_data = 12'b110011001001;
		if(({row_reg, col_reg}==16'b0010111100011101)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==16'b0010111100011110)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0010111100011111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0010111100100000) && ({row_reg, col_reg}<16'b0010111100100101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010111100100101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0010111100100110)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0010111100100111)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0010111100101000)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0010111100101001)) color_data = 12'b110011001001;
		if(({row_reg, col_reg}==16'b0010111100101010)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0010111100101011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0010111100101100)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=16'b0010111100101101) && ({row_reg, col_reg}<16'b0010111100101111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010111100101111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0010111100110000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0010111100110001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0010111100110010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0010111100110011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010111100110100)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0010111100110101)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==16'b0010111100110110)) color_data = 12'b100010010111;
		if(({row_reg, col_reg}>=16'b0010111100110111) && ({row_reg, col_reg}<16'b0010111100111001)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0010111100111001)) color_data = 12'b100110101000;
		if(({row_reg, col_reg}==16'b0010111100111010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0010111100111011)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0010111100111100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0010111100111101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0010111100111110) && ({row_reg, col_reg}<16'b0010111101000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010111101000000) && ({row_reg, col_reg}<16'b0010111101000010)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0010111101000010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010111101000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111101000100) && ({row_reg, col_reg}<16'b0010111101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111101000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010111101000111) && ({row_reg, col_reg}<16'b0010111101001001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010111101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111101001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010111101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111101001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010111101001110) && ({row_reg, col_reg}<16'b0010111101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111101010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010111101010001) && ({row_reg, col_reg}<16'b0010111101010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010111101010011) && ({row_reg, col_reg}<16'b0010111101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010111101011110) && ({row_reg, col_reg}<16'b0010111101100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111101100000) && ({row_reg, col_reg}<16'b0010111101100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111101100011) && ({row_reg, col_reg}<16'b0010111101100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111101100101) && ({row_reg, col_reg}<16'b0010111101100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010111101100111) && ({row_reg, col_reg}<16'b0010111101101001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010111101101001) && ({row_reg, col_reg}<16'b0010111101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111101101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010111101101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111101101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010111101101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111101110000) && ({row_reg, col_reg}<16'b0010111101110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111101110010) && ({row_reg, col_reg}<16'b0010111101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010111101110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010111101110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010111101110110) && ({row_reg, col_reg}<16'b0010111101111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010111101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111101111001) && ({row_reg, col_reg}<16'b0010111101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111101111100) && ({row_reg, col_reg}<16'b0010111101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010111101111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010111110000000) && ({row_reg, col_reg}<16'b0010111110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111110000011) && ({row_reg, col_reg}<16'b0010111110100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010111110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111110100101) && ({row_reg, col_reg}<16'b0010111110101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111110101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111110101001) && ({row_reg, col_reg}<16'b0010111110101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010111110101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111110110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111110110001) && ({row_reg, col_reg}<16'b0010111110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010111110110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111110110100) && ({row_reg, col_reg}<16'b0010111110110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111110110110) && ({row_reg, col_reg}<16'b0010111110111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111110111000) && ({row_reg, col_reg}<16'b0010111110111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111110111010) && ({row_reg, col_reg}<16'b0010111111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111111000000) && ({row_reg, col_reg}<16'b0010111111000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111111000101) && ({row_reg, col_reg}<16'b0010111111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111111001001) && ({row_reg, col_reg}<16'b0010111111001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111111001011) && ({row_reg, col_reg}<16'b0010111111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111111001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111111001111) && ({row_reg, col_reg}<16'b0010111111010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111111010010) && ({row_reg, col_reg}<16'b0010111111010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111111010100) && ({row_reg, col_reg}<16'b0010111111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111111011111) && ({row_reg, col_reg}<16'b0010111111100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111111100010) && ({row_reg, col_reg}<16'b0010111111100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111111100101) && ({row_reg, col_reg}<16'b0010111111100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111111100111) && ({row_reg, col_reg}<16'b0010111111101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111111101010) && ({row_reg, col_reg}<16'b0010111111101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010111111101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111111101110) && ({row_reg, col_reg}<16'b0010111111110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111111110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111111110001)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0010111111110010) && ({row_reg, col_reg}<16'b0011000000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011000000000000) && ({row_reg, col_reg}<16'b0011000000000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000000000010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0011000000000011) && ({row_reg, col_reg}<16'b0011000000000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011000000000101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0011000000000110) && ({row_reg, col_reg}<16'b0011000000001001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011000000001001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011000000001010)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011000000001011)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==16'b0011000000001100)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011000000001101)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==16'b0011000000001110)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011000000001111)) color_data = 12'b100110101000;
		if(({row_reg, col_reg}==16'b0011000000010000)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011000000010001)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=16'b0011000000010010) && ({row_reg, col_reg}<16'b0011000000010101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011000000010101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011000000010110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011000000010111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011000000011000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011000000011001)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==16'b0011000000011010)) color_data = 12'b101010111001;
		if(({row_reg, col_reg}==16'b0011000000011011)) color_data = 12'b110011011010;
		if(({row_reg, col_reg}==16'b0011000000011100)) color_data = 12'b101111001001;
		if(({row_reg, col_reg}==16'b0011000000011101)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011000000011110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0011000000011111) && ({row_reg, col_reg}<16'b0011000000100001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011000000100001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0011000000100010) && ({row_reg, col_reg}<16'b0011000000100101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011000000100101)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011000000100110)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011000000100111)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011000000101000)) color_data = 12'b110111011010;
		if(({row_reg, col_reg}==16'b0011000000101001)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==16'b0011000000101010)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011000000101011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011000000101100)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011000000101101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011000000101110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011000000101111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011000000110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011000000110001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011000000110010)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011000000110011)) color_data = 12'b100010010111;
		if(({row_reg, col_reg}>=16'b0011000000110100) && ({row_reg, col_reg}<16'b0011000000110110)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011000000110110)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011000000110111)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011000000111000)) color_data = 12'b100110101000;
		if(({row_reg, col_reg}==16'b0011000000111001)) color_data = 12'b011110000110;
		if(({row_reg, col_reg}==16'b0011000000111010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011000000111011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011000000111100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011000000111101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011000000111110)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0011000000111111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011000001000000) && ({row_reg, col_reg}<16'b0011000001000010)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0011000001000010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011000001000011) && ({row_reg, col_reg}<16'b0011000001000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000001000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011000001000111) && ({row_reg, col_reg}<16'b0011000001001001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011000001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000001001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011000001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011000001001100) && ({row_reg, col_reg}<16'b0011000001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000001010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011000001010001) && ({row_reg, col_reg}<16'b0011000001010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011000001010011) && ({row_reg, col_reg}<16'b0011000001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000001011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011000001100000) && ({row_reg, col_reg}<16'b0011000001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000001100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011000001100011) && ({row_reg, col_reg}<16'b0011000001100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011000001100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011000001100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000001100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011000001101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011000001101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000001101010) && ({row_reg, col_reg}<16'b0011000001101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000001101100) && ({row_reg, col_reg}<16'b0011000001101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000001101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011000001101111) && ({row_reg, col_reg}<16'b0011000001110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000001110010) && ({row_reg, col_reg}<16'b0011000001110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011000001110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000001110101) && ({row_reg, col_reg}<16'b0011000001110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011000001110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000001111000) && ({row_reg, col_reg}<16'b0011000001111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000001111010) && ({row_reg, col_reg}<16'b0011000001111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011000001111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000001111101) && ({row_reg, col_reg}<16'b0011000010000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011000010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011000010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000010000011) && ({row_reg, col_reg}<16'b0011000010100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011000010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000010100101) && ({row_reg, col_reg}<16'b0011000010101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011000010101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000010101001) && ({row_reg, col_reg}<16'b0011000010101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011000010101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000010110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000010110001) && ({row_reg, col_reg}<16'b0011000010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011000010110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000010110100) && ({row_reg, col_reg}<16'b0011000010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000010110110) && ({row_reg, col_reg}<16'b0011000010111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000010111100) && ({row_reg, col_reg}<16'b0011000010111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000010111110) && ({row_reg, col_reg}<16'b0011000011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000011000000) && ({row_reg, col_reg}<16'b0011000011000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000011000011) && ({row_reg, col_reg}<16'b0011000011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000011001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000011001010) && ({row_reg, col_reg}<16'b0011000011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000011001110) && ({row_reg, col_reg}<16'b0011000011010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000011010100) && ({row_reg, col_reg}<16'b0011000011010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000011010110) && ({row_reg, col_reg}<16'b0011000011011011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011000011011011) && ({row_reg, col_reg}<16'b0011000011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000011011111) && ({row_reg, col_reg}<16'b0011000011100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000011100011) && ({row_reg, col_reg}<16'b0011000011100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000011100101) && ({row_reg, col_reg}<16'b0011000011101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011000011101100) && ({row_reg, col_reg}<16'b0011000011101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000011101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000011101111) && ({row_reg, col_reg}<16'b0011000011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000011110001)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0011000011110010) && ({row_reg, col_reg}<16'b0011000100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011000100000000) && ({row_reg, col_reg}<16'b0011000100000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000100000011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011000100000100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011000100000101) && ({row_reg, col_reg}<16'b0011000100000111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0011000100000111) && ({row_reg, col_reg}<16'b0011000100001010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011000100001010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011000100001011)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011000100001100)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==16'b0011000100001101)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011000100001110)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==16'b0011000100001111)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011000100010000)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011000100010001)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011000100010010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011000100010011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0011000100010100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011000100010101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011000100010110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011000100010111)) color_data = 12'b010101100100;
		if(({row_reg, col_reg}==16'b0011000100011000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011000100011001)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011000100011010)) color_data = 12'b110011001001;
		if(({row_reg, col_reg}==16'b0011000100011011)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==16'b0011000100011100)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011000100011101)) color_data = 12'b010101100100;
		if(({row_reg, col_reg}==16'b0011000100011110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011000100011111) && ({row_reg, col_reg}<16'b0011000100100011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011000100100011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011000100100100)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011000100100101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011000100100110)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}>=16'b0011000100100111) && ({row_reg, col_reg}<16'b0011000100101001)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011000100101001)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011000100101010)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011000100101011)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011000100101100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011000100101101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0011000100101110) && ({row_reg, col_reg}<16'b0011000100110000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011000100110000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011000100110001)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011000100110010)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011000100110011)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011000100110100)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011000100110101)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}>=16'b0011000100110110) && ({row_reg, col_reg}<16'b0011000100111000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011000100111000)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011000100111001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011000100111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011000100111011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011000100111100)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011000100111101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011000100111110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011000100111111) && ({row_reg, col_reg}<16'b0011000101000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011000101000011) && ({row_reg, col_reg}<16'b0011000101000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000101000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011000101000111) && ({row_reg, col_reg}<16'b0011000101001001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011000101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011000101001010) && ({row_reg, col_reg}<16'b0011000101001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000101001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011000101001110) && ({row_reg, col_reg}<16'b0011000101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000101010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011000101010001) && ({row_reg, col_reg}<16'b0011000101010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011000101010011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011000101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000101010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011000101010110) && ({row_reg, col_reg}<16'b0011000101011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011000101011000) && ({row_reg, col_reg}<16'b0011000101011010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011000101011010) && ({row_reg, col_reg}<16'b0011000101100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011000101100011) && ({row_reg, col_reg}<16'b0011000101100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011000101100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011000101100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000101100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011000101101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011000101101001) && ({row_reg, col_reg}<16'b0011000101101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000101101011) && ({row_reg, col_reg}<16'b0011000101101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011000101101110) && ({row_reg, col_reg}<16'b0011000101110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000101110000) && ({row_reg, col_reg}<16'b0011000101110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000101110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011000101110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011000101110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011000101110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011000101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000101110111) && ({row_reg, col_reg}<16'b0011000101111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000101111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011000101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000101111100) && ({row_reg, col_reg}<16'b0011000101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000101111110) && ({row_reg, col_reg}<16'b0011000110000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011000110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011000110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000110000011) && ({row_reg, col_reg}<16'b0011000110100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011000110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000110100101) && ({row_reg, col_reg}<16'b0011000110100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000110100111) && ({row_reg, col_reg}<16'b0011000110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000110101001) && ({row_reg, col_reg}<16'b0011000110101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011000110101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000110110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000110110001) && ({row_reg, col_reg}<16'b0011000110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011000110110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000110110100) && ({row_reg, col_reg}<16'b0011000110111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000110111010) && ({row_reg, col_reg}<16'b0011000110111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000110111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000110111101) && ({row_reg, col_reg}<16'b0011000111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000111000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000111000010) && ({row_reg, col_reg}<16'b0011000111001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000111001101) && ({row_reg, col_reg}<16'b0011000111010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011000111010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000111010110) && ({row_reg, col_reg}<16'b0011000111011000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011000111011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000111011001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011000111011010) && ({row_reg, col_reg}<16'b0011000111011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000111011110) && ({row_reg, col_reg}<16'b0011000111100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000111100011) && ({row_reg, col_reg}<16'b0011000111100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000111100111) && ({row_reg, col_reg}<16'b0011000111101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011000111101010) && ({row_reg, col_reg}<16'b0011000111110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000111110000) && ({row_reg, col_reg}<16'b0011000111110010)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0011000111110010) && ({row_reg, col_reg}<16'b0011001000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011001000000000) && ({row_reg, col_reg}<16'b0011001000000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001000000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011001000000100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011001000000101)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011001000000110)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011001000000111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0011001000001000) && ({row_reg, col_reg}<16'b0011001000001011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011001000001011)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011001000001100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011001000001101)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011001000001110)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==16'b0011001000001111)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011001000010000)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011001000010001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0011001000010010) && ({row_reg, col_reg}<16'b0011001000010101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011001000010101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011001000010110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011001000010111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011001000011000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011001000011001)) color_data = 12'b101110111000;
		if(({row_reg, col_reg}==16'b0011001000011010)) color_data = 12'b110011001001;
		if(({row_reg, col_reg}==16'b0011001000011011)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011001000011100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011001000011101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011001000011110)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}>=16'b0011001000011111) && ({row_reg, col_reg}<16'b0011001000100001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011001000100001)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0011001000100010)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0011001000100011)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011001000100100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011001000100101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011001000100110)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==16'b0011001000100111)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011001000101000)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==16'b0011001000101001)) color_data = 12'b100001110101;
		if(({row_reg, col_reg}==16'b0011001000101010)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0011001000101011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011001000101100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0011001000101101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011001000101110)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}>=16'b0011001000101111) && ({row_reg, col_reg}<16'b0011001000110001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011001000110001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011001000110010)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011001000110011)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==16'b0011001000110100)) color_data = 12'b100001110101;
		if(({row_reg, col_reg}==16'b0011001000110101)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}>=16'b0011001000110110) && ({row_reg, col_reg}<16'b0011001000111010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011001000111010)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}>=16'b0011001000111011) && ({row_reg, col_reg}<16'b0011001000111101)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011001000111101)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==16'b0011001000111110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0011001000111111) && ({row_reg, col_reg}<16'b0011001001000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011001001000011) && ({row_reg, col_reg}<16'b0011001001000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011001001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001001000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011001001000111) && ({row_reg, col_reg}<16'b0011001001001001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011001001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011001001001010) && ({row_reg, col_reg}<16'b0011001001001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001001001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001001001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011001001001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001001010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011001001010001) && ({row_reg, col_reg}<16'b0011001001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011001001010100) && ({row_reg, col_reg}<16'b0011001001011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011001001011000) && ({row_reg, col_reg}<16'b0011001001011011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011001001011011) && ({row_reg, col_reg}<16'b0011001001011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001001011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011001001011110) && ({row_reg, col_reg}<16'b0011001001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001001100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011001001100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011001001100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001001100101) && ({row_reg, col_reg}<16'b0011001001100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011001001100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011001001101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011001001101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001001101010) && ({row_reg, col_reg}<16'b0011001001101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011001001101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011001001101101) && ({row_reg, col_reg}<16'b0011001001110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011001001110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011001001110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001001110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011001001110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011001001110100) && ({row_reg, col_reg}<16'b0011001001110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001001110110) && ({row_reg, col_reg}<16'b0011001001111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001001111001) && ({row_reg, col_reg}<16'b0011001001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011001001111011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=16'b0011001001111100) && ({row_reg, col_reg}<16'b0011001001111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011001001111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011001010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011001010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001010000011) && ({row_reg, col_reg}<16'b0011001010100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011001010100100) && ({row_reg, col_reg}<16'b0011001010100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001010100111) && ({row_reg, col_reg}<16'b0011001010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001010101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011001010101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011001010101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011001010101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011001010101110) && ({row_reg, col_reg}<16'b0011001010110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001010110001) && ({row_reg, col_reg}<16'b0011001010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011001010110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001010110100) && ({row_reg, col_reg}<16'b0011001010111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001010111010) && ({row_reg, col_reg}<16'b0011001010111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001010111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001010111101) && ({row_reg, col_reg}<16'b0011001011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001011000010) && ({row_reg, col_reg}<16'b0011001011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001011001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001011001010) && ({row_reg, col_reg}<16'b0011001011001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001011001101) && ({row_reg, col_reg}<16'b0011001011001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001011001111) && ({row_reg, col_reg}<16'b0011001011010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001011010010) && ({row_reg, col_reg}<16'b0011001011010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001011010110) && ({row_reg, col_reg}<16'b0011001011011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001011011101) && ({row_reg, col_reg}<16'b0011001011100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001011100001) && ({row_reg, col_reg}<16'b0011001011101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001011101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011001011101001) && ({row_reg, col_reg}<16'b0011001011110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001011110000)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0011001011110001) && ({row_reg, col_reg}<16'b0011001100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011001100000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011001100000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001100000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011001100000011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011001100000100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011001100000101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011001100000110)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==16'b0011001100000111)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011001100001000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011001100001001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011001100001010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011001100001011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011001100001100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011001100001101)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011001100001110)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011001100001111)) color_data = 12'b101110101000;
		if(({row_reg, col_reg}==16'b0011001100010000)) color_data = 12'b100001110101;
		if(({row_reg, col_reg}>=16'b0011001100010001) && ({row_reg, col_reg}<16'b0011001100010101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011001100010101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011001100010110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011001100010111)) color_data = 12'b010101100100;
		if(({row_reg, col_reg}==16'b0011001100011000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011001100011001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==16'b0011001100011010)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011001100011011)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011001100011100)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011001100011101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0011001100011110) && ({row_reg, col_reg}<16'b0011001100100000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011001100100000) && ({row_reg, col_reg}<16'b0011001100100010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011001100100010)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011001100100011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011001100100100)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==16'b0011001100100101)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}>=16'b0011001100100110) && ({row_reg, col_reg}<16'b0011001100101000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011001100101000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011001100101001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011001100101010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0011001100101011) && ({row_reg, col_reg}<16'b0011001100101101)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0011001100101101)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011001100101110)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==16'b0011001100101111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=16'b0011001100110000) && ({row_reg, col_reg}<16'b0011001100110010)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011001100110010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011001100110011)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011001100110100)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011001100110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011001100110110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011001100110111)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0011001100111000)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0011001100111001)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011001100111010)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011001100111011)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011001100111100)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==16'b0011001100111101)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011001100111110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011001100111111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011001101000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011001101000001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0011001101000010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011001101000011) && ({row_reg, col_reg}<16'b0011001101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001101000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011001101000111) && ({row_reg, col_reg}<16'b0011001101001001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011001101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011001101001010) && ({row_reg, col_reg}<16'b0011001101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001101001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011001101001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001101001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011001101001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001101010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011001101010001) && ({row_reg, col_reg}<16'b0011001101010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011001101010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011001101010100) && ({row_reg, col_reg}<16'b0011001101010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001101010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011001101010111) && ({row_reg, col_reg}<16'b0011001101011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011001101011001) && ({row_reg, col_reg}<16'b0011001101011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011001101011110) && ({row_reg, col_reg}<16'b0011001101100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001101100010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011001101100011) && ({row_reg, col_reg}<16'b0011001101100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001101100101) && ({row_reg, col_reg}<16'b0011001101100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011001101100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011001101101000) && ({row_reg, col_reg}<16'b0011001101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001101101010) && ({row_reg, col_reg}<16'b0011001101101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011001101101100) && ({row_reg, col_reg}<16'b0011001101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001101101110) && ({row_reg, col_reg}<16'b0011001101110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011001101110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011001101110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001101110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011001101110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011001101110100) && ({row_reg, col_reg}<16'b0011001101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001101110110) && ({row_reg, col_reg}<16'b0011001101111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001101111001) && ({row_reg, col_reg}<16'b0011001101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011001101111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011001101111100) && ({row_reg, col_reg}<16'b0011001101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001101111111) && ({row_reg, col_reg}<16'b0011001110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011001110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001110000011) && ({row_reg, col_reg}<16'b0011001110100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011001110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001110100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011001110100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001110100111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001110101000) && ({row_reg, col_reg}<16'b0011001110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001110101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011001110101011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==16'b0011001110101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001110101101) && ({row_reg, col_reg}<16'b0011001110110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001110110000) && ({row_reg, col_reg}<16'b0011001110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011001110110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001110110100) && ({row_reg, col_reg}<16'b0011001110111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001110111010) && ({row_reg, col_reg}<16'b0011001110111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001110111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001110111101) && ({row_reg, col_reg}<16'b0011001111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001111001001) && ({row_reg, col_reg}<16'b0011001111001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001111001011) && ({row_reg, col_reg}<16'b0011001111001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001111001101) && ({row_reg, col_reg}<16'b0011001111001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001111001111) && ({row_reg, col_reg}<16'b0011001111010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001111010010) && ({row_reg, col_reg}<16'b0011001111010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001111010110) && ({row_reg, col_reg}<16'b0011001111011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001111011101) && ({row_reg, col_reg}<16'b0011001111011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001111011111) && ({row_reg, col_reg}<16'b0011001111100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001111100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001111100011) && ({row_reg, col_reg}<16'b0011001111110000)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0011001111110000) && ({row_reg, col_reg}<16'b0011010000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011010000000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010000000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010000000010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0011010000000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010000000100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011010000000101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011010000000110)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==16'b0011010000000111)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011010000001000)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0011010000001001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011010000001010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011010000001011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011010000001100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011010000001101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011010000001110)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011010000001111)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==16'b0011010000010000)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==16'b0011010000010001)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011010000010010)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0011010000010011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011010000010100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0011010000010101) && ({row_reg, col_reg}<16'b0011010000010111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011010000010111)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011010000011000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011010000011001)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==16'b0011010000011010)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011010000011011)) color_data = 12'b100001110101;
		if(({row_reg, col_reg}==16'b0011010000011100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0011010000011101) && ({row_reg, col_reg}<16'b0011010000011111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011010000011111)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011010000100000)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011010000100001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011010000100010)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011010000100011)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011010000100100)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011010000100101)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0011010000100110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011010000100111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0011010000101000) && ({row_reg, col_reg}<16'b0011010000101010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011010000101010)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011010000101011)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011010000101100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011010000101101)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==16'b0011010000101110)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011010000101111)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0011010000110000)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011010000110001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011010000110010)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0011010000110011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011010000110100)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011010000110101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011010000110110)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011010000110111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011010000111000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011010000111001)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011010000111010)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011010000111011)) color_data = 12'b110011001001;
		if(({row_reg, col_reg}==16'b0011010000111100)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==16'b0011010000111101)) color_data = 12'b110011011010;
		if(({row_reg, col_reg}==16'b0011010000111110)) color_data = 12'b100110101000;
		if(({row_reg, col_reg}==16'b0011010000111111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011010001000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011010001000001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011010001000010)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0011010001000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011010001000100) && ({row_reg, col_reg}<16'b0011010001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010001000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011010001000111) && ({row_reg, col_reg}<16'b0011010001001001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011010001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011010001001010) && ({row_reg, col_reg}<16'b0011010001001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010001001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011010001001110) && ({row_reg, col_reg}<16'b0011010001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010001010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011010001010001) && ({row_reg, col_reg}<16'b0011010001010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011010001010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011010001010100) && ({row_reg, col_reg}<16'b0011010001010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010001010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011010001010111) && ({row_reg, col_reg}<16'b0011010001011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011010001011001) && ({row_reg, col_reg}<16'b0011010001011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011010001011110) && ({row_reg, col_reg}<16'b0011010001100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011010001100001) && ({row_reg, col_reg}<16'b0011010001100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011010001100011) && ({row_reg, col_reg}<16'b0011010001100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011010001100101) && ({row_reg, col_reg}<16'b0011010001100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011010001100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011010001101000) && ({row_reg, col_reg}<16'b0011010001101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011010001101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010001101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011010001101100) && ({row_reg, col_reg}<16'b0011010001101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010001101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011010001101111) && ({row_reg, col_reg}<16'b0011010001110001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011010001110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010001110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011010001110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011010001110100) && ({row_reg, col_reg}<16'b0011010001110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010001110110) && ({row_reg, col_reg}<16'b0011010001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010001111000) && ({row_reg, col_reg}<16'b0011010001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010001111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011010001111100) && ({row_reg, col_reg}<16'b0011010010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010010000000) && ({row_reg, col_reg}<16'b0011010010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010010000011) && ({row_reg, col_reg}<16'b0011010010100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011010010100100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010010100101) && ({row_reg, col_reg}<16'b0011010010100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010010100111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010010101000) && ({row_reg, col_reg}<16'b0011010010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010010101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010010101011) && ({row_reg, col_reg}<16'b0011010010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011010010110000) && ({row_reg, col_reg}<16'b0011010010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011010010110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010010110100) && ({row_reg, col_reg}<16'b0011010010111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011010010111001) && ({row_reg, col_reg}<16'b0011010011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010011001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010011001011) && ({row_reg, col_reg}<16'b0011010011001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010011001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010011001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011010011001111) && ({row_reg, col_reg}<16'b0011010011010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010011010001) && ({row_reg, col_reg}<16'b0011010011011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010011011101)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==16'b0011010011011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011010011011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011010011100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010011100001) && ({row_reg, col_reg}<16'b0011010011100110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010011100110) && ({row_reg, col_reg}<16'b0011010011101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010011101011) && ({row_reg, col_reg}<16'b0011010011101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010011101110) && ({row_reg, col_reg}<16'b0011010011110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010011110000)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0011010011110001) && ({row_reg, col_reg}<16'b0011010100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011010100000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010100000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010100000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010100000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010100000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011010100000101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011010100000110)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011010100000111)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011010100001000)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=16'b0011010100001001) && ({row_reg, col_reg}<16'b0011010100001011)) color_data = 12'b100001110101;
		if(({row_reg, col_reg}==16'b0011010100001011)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011010100001100)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011010100001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011010100001110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0011010100001111) && ({row_reg, col_reg}<16'b0011010100010001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011010100010001)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011010100010010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0011010100010011) && ({row_reg, col_reg}<16'b0011010100010111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011010100010111)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}>=16'b0011010100011000) && ({row_reg, col_reg}<16'b0011010100011010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011010100011010)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011010100011011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011010100011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0011010100011101) && ({row_reg, col_reg}<16'b0011010100011111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011010100011111)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011010100100000)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011010100100001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011010100100010)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011010100100011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011010100100100)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011010100100101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011010100100110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011010100100111) && ({row_reg, col_reg}<16'b0011010100101001)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0011010100101001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011010100101010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=16'b0011010100101011) && ({row_reg, col_reg}<16'b0011010100101101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011010100101101)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011010100101110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0011010100101111) && ({row_reg, col_reg}<16'b0011010100110001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0011010100110001) && ({row_reg, col_reg}<16'b0011010100110011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011010100110011)) color_data = 12'b011001110101;
		if(({row_reg, col_reg}==16'b0011010100110100)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==16'b0011010100110101)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011010100110110)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==16'b0011010100110111)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0011010100111000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011010100111001)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011010100111010)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==16'b0011010100111011)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}>=16'b0011010100111100) && ({row_reg, col_reg}<16'b0011010100111110)) color_data = 12'b101110111000;
		if(({row_reg, col_reg}==16'b0011010100111110)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011010100111111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011010101000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011010101000001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0011010101000010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011010101000011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011010101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010101000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011010101000111) && ({row_reg, col_reg}<16'b0011010101001001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011010101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011010101001010) && ({row_reg, col_reg}<16'b0011010101001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010101001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011010101001110) && ({row_reg, col_reg}<16'b0011010101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011010101010000) && ({row_reg, col_reg}<16'b0011010101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011010101010100) && ({row_reg, col_reg}<16'b0011010101010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010101010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011010101010111) && ({row_reg, col_reg}<16'b0011010101011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011010101011001) && ({row_reg, col_reg}<16'b0011010101011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011010101011110) && ({row_reg, col_reg}<16'b0011010101100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011010101100011) && ({row_reg, col_reg}<16'b0011010101100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011010101100101) && ({row_reg, col_reg}<16'b0011010101100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011010101100111) && ({row_reg, col_reg}<16'b0011010101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010101101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011010101101011) && ({row_reg, col_reg}<16'b0011010101110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010101110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010101110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011010101110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011010101110100) && ({row_reg, col_reg}<16'b0011010101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010101110110) && ({row_reg, col_reg}<16'b0011010101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010101111000) && ({row_reg, col_reg}<16'b0011010101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010101111100) && ({row_reg, col_reg}<16'b0011010110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010110000000) && ({row_reg, col_reg}<16'b0011010110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010110000011) && ({row_reg, col_reg}<16'b0011010110100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011010110100100) && ({row_reg, col_reg}<16'b0011010110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010110101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011010110101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011010110101011) && ({row_reg, col_reg}<16'b0011010110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011010110110000) && ({row_reg, col_reg}<16'b0011010110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011010110110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010110110100) && ({row_reg, col_reg}<16'b0011010110110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011010110110111) && ({row_reg, col_reg}<16'b0011010110111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010110111010) && ({row_reg, col_reg}<16'b0011010110111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010110111100) && ({row_reg, col_reg}<16'b0011010110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010110111110) && ({row_reg, col_reg}<16'b0011010111000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010111000001) && ({row_reg, col_reg}<16'b0011010111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010111000111) && ({row_reg, col_reg}<16'b0011010111001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010111001001) && ({row_reg, col_reg}<16'b0011010111001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010111001101) && ({row_reg, col_reg}<16'b0011010111001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011010111001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011010111010000) && ({row_reg, col_reg}<16'b0011010111010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010111010010) && ({row_reg, col_reg}<16'b0011010111010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010111010101) && ({row_reg, col_reg}<16'b0011010111011110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011010111011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011010111011111) && ({row_reg, col_reg}<16'b0011010111100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011010111100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010111100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011010111100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011010111100100) && ({row_reg, col_reg}<16'b0011010111100110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010111100110) && ({row_reg, col_reg}<16'b0011010111110001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0011010111110001) && ({row_reg, col_reg}<16'b0011011000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011011000000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011011000000001) && ({row_reg, col_reg}<16'b0011011000000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011000000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011011000000100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011011000000101) && ({row_reg, col_reg}<16'b0011011000001000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011011000001000)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==16'b0011011000001001)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011011000001010)) color_data = 12'b110011001001;
		if(({row_reg, col_reg}==16'b0011011000001011)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011011000001100)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011011000001101)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0011011000001110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011011000001111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011011000010000)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}>=16'b0011011000010001) && ({row_reg, col_reg}<16'b0011011000010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011011000010100) && ({row_reg, col_reg}<16'b0011011000010111)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0011011000010111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011011000011000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011011000011001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0011011000011010)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0011011000011011) && ({row_reg, col_reg}<16'b0011011000011110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011011000011110) && ({row_reg, col_reg}<16'b0011011000100000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011011000100000) && ({row_reg, col_reg}<16'b0011011000100101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011011000100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011011000100110)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0011011000100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011011000101000)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0011011000101001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0011011000101010) && ({row_reg, col_reg}<16'b0011011000101100)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0011011000101100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0011011000101101) && ({row_reg, col_reg}<16'b0011011000101111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0011011000101111) && ({row_reg, col_reg}<16'b0011011000110001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011011000110001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011011000110010)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011011000110011)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011011000110100)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011011000110101)) color_data = 12'b110111011010;
		if(({row_reg, col_reg}==16'b0011011000110110)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011011000110111)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011011000111000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011011000111001)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011011000111010)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==16'b0011011000111011)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011011000111100)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011011000111101)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011011000111110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011011000111111)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0011011001000000) && ({row_reg, col_reg}<16'b0011011001000010)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0011011001000010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011011001000011) && ({row_reg, col_reg}<16'b0011011001000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011001000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011011001000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011011001001000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011011001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011011001001010) && ({row_reg, col_reg}<16'b0011011001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011001001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011011001001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011011001001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011011001001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011011001010000) && ({row_reg, col_reg}<16'b0011011001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011011001010100) && ({row_reg, col_reg}<16'b0011011001010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011001010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011011001010111) && ({row_reg, col_reg}<16'b0011011001011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011011001011001) && ({row_reg, col_reg}<16'b0011011001011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011011001011110) && ({row_reg, col_reg}<16'b0011011001100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011011001100001) && ({row_reg, col_reg}<16'b0011011001100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011011001100011) && ({row_reg, col_reg}<16'b0011011001100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011011001100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011011001100110) && ({row_reg, col_reg}<16'b0011011001101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011011001101001) && ({row_reg, col_reg}<16'b0011011001101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011011001101100) && ({row_reg, col_reg}<16'b0011011001110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011001110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011001110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011011001110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011011001110100) && ({row_reg, col_reg}<16'b0011011001110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011001110110) && ({row_reg, col_reg}<16'b0011011001111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011001111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011001111010) && ({row_reg, col_reg}<16'b0011011010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011010000010) && ({row_reg, col_reg}<16'b0011011010100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011011010100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011010100101) && ({row_reg, col_reg}<16'b0011011010101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011010101001) && ({row_reg, col_reg}<16'b0011011010101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011010101011) && ({row_reg, col_reg}<16'b0011011010101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011010101110) && ({row_reg, col_reg}<16'b0011011010110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011010110000) && ({row_reg, col_reg}<16'b0011011010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011011010110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011010110100) && ({row_reg, col_reg}<16'b0011011010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011010110111) && ({row_reg, col_reg}<16'b0011011010111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011011010111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011010111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011010111100) && ({row_reg, col_reg}<16'b0011011010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011010111110) && ({row_reg, col_reg}<16'b0011011011000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011011000000) && ({row_reg, col_reg}<16'b0011011011000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011011011000010) && ({row_reg, col_reg}<16'b0011011011000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011011000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011011011000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011011000111) && ({row_reg, col_reg}<16'b0011011011001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011011001001) && ({row_reg, col_reg}<16'b0011011011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011011001110) && ({row_reg, col_reg}<16'b0011011011010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011011011010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011011010011) && ({row_reg, col_reg}<16'b0011011011011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011011011011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011011011101) && ({row_reg, col_reg}<16'b0011011011100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011011011100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011011100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011011100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011011100100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011011100101) && ({row_reg, col_reg}<16'b0011011011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011011101111) && ({row_reg, col_reg}<16'b0011011011110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011011110001) && ({row_reg, col_reg}<16'b0011011011111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011011011111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0011011011111100) && ({row_reg, col_reg}<16'b0011011100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011011100000000) && ({row_reg, col_reg}<16'b0011011100000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011100000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011011100000100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011011100000101) && ({row_reg, col_reg}<16'b0011011100001000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011011100001000)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011011100001001)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011011100001010)) color_data = 12'b110111101011;
		if(({row_reg, col_reg}==16'b0011011100001011)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==16'b0011011100001100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011011100001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011011100001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011100010000) && ({row_reg, col_reg}<16'b0011011100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011100010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011011100010100) && ({row_reg, col_reg}<16'b0011011100011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011011100011001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011011100011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011100011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011011100011100) && ({row_reg, col_reg}<16'b0011011100011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011011100011111)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0011011100100000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011011100100001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0011011100100010) && ({row_reg, col_reg}<16'b0011011100100100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011011100100100) && ({row_reg, col_reg}<16'b0011011100100110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011011100100110)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0011011100100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011011100101000)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0011011100101001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011011100101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011011100101011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011011100101100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0011011100101101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0011011100101110)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}>=16'b0011011100101111) && ({row_reg, col_reg}<16'b0011011100110001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011011100110001)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0011011100110010)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011011100110011)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011011100110100)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011011100110101)) color_data = 12'b101110111000;
		if(({row_reg, col_reg}==16'b0011011100110110)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011011100110111)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0011011100111000)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0011011100111001)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011011100111010)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011011100111011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011011100111100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0011011100111101) && ({row_reg, col_reg}<16'b0011011101000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011011101000000)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0011011101000001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0011011101000010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011011101000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011101000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011011101000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011011101001000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011011101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011011101001010) && ({row_reg, col_reg}<16'b0011011101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011011101001100) && ({row_reg, col_reg}<16'b0011011101001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011011101001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011011101001111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0011011101010000) && ({row_reg, col_reg}<16'b0011011101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011011101010100) && ({row_reg, col_reg}<16'b0011011101011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011011101011011) && ({row_reg, col_reg}<16'b0011011101011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011011101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011011101011111) && ({row_reg, col_reg}<16'b0011011101100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011011101100011) && ({row_reg, col_reg}<16'b0011011101100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011011101100101) && ({row_reg, col_reg}<16'b0011011101100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011011101100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011011101101000) && ({row_reg, col_reg}<16'b0011011101101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011011101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011101101101) && ({row_reg, col_reg}<16'b0011011101101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011011101101111) && ({row_reg, col_reg}<16'b0011011101110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011101110010) && ({row_reg, col_reg}<16'b0011011101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011011101110100) && ({row_reg, col_reg}<16'b0011011101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011101110110) && ({row_reg, col_reg}<16'b0011011101111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011101111001) && ({row_reg, col_reg}<16'b0011011101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011101111011) && ({row_reg, col_reg}<16'b0011011110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011110000010) && ({row_reg, col_reg}<16'b0011011110100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011011110100100) && ({row_reg, col_reg}<16'b0011011110100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011110100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011110100111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011110101000) && ({row_reg, col_reg}<16'b0011011110101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011110101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011110101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011011110101111) && ({row_reg, col_reg}<16'b0011011110110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011110110001) && ({row_reg, col_reg}<16'b0011011110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011011110110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011110110100) && ({row_reg, col_reg}<16'b0011011110110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011110110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011011110110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011011110111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011110111001) && ({row_reg, col_reg}<16'b0011011110111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011110111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011111000000) && ({row_reg, col_reg}<16'b0011011111000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011011111000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011111000011) && ({row_reg, col_reg}<16'b0011011111011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011111011110) && ({row_reg, col_reg}<16'b0011011111100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011011111100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011111100010) && ({row_reg, col_reg}<16'b0011011111100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011111100100) && ({row_reg, col_reg}<16'b0011011111100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011111100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011011111101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011111101001) && ({row_reg, col_reg}<16'b0011011111101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011011111101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011111101101) && ({row_reg, col_reg}<16'b0011011111101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011011111101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011111110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011111110001) && ({row_reg, col_reg}<16'b0011011111111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011011111111010) && ({row_reg, col_reg}<16'b0011011111111100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0011011111111100) && ({row_reg, col_reg}<16'b0011100000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011100000000000) && ({row_reg, col_reg}<16'b0011100000000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100000000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011100000000100) && ({row_reg, col_reg}<16'b0011100000001000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011100000001000)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011100000001001)) color_data = 12'b100010010111;
		if(({row_reg, col_reg}>=16'b0011100000001010) && ({row_reg, col_reg}<16'b0011100000001100)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011100000001100)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011100000001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011100000001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011100000001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100000010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011100000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011100000010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100000010011) && ({row_reg, col_reg}<16'b0011100000010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011100000010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100000010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100000010111) && ({row_reg, col_reg}<16'b0011100000011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100000011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100000011010) && ({row_reg, col_reg}<16'b0011100000011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011100000011100) && ({row_reg, col_reg}<16'b0011100000101111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011100000101111)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0011100000110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011100000110001)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011100000110010)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011100000110011)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011100000110100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011100000110101)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011100000110110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011100000110111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011100000111000)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0011100000111001) && ({row_reg, col_reg}<16'b0011100000111011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011100000111011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0011100000111100) && ({row_reg, col_reg}<16'b0011100001000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011100001000000)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0011100001000001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0011100001000010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011100001000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011100001000100) && ({row_reg, col_reg}<16'b0011100001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100001000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011100001000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011100001001000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011100001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011100001001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011100001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011100001001100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011100001001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011100001001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011100001001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011100001010000) && ({row_reg, col_reg}<16'b0011100001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011100001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100001010101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0011100001010110) && ({row_reg, col_reg}<16'b0011100001011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011100001011000) && ({row_reg, col_reg}<16'b0011100001011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011100001011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100001011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011100001100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011100001100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011100001100010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011100001100011) && ({row_reg, col_reg}<16'b0011100001100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100001100101) && ({row_reg, col_reg}<16'b0011100001101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011100001101100) && ({row_reg, col_reg}<16'b0011100001101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011100001101110) && ({row_reg, col_reg}<16'b0011100001110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011100001110000) && ({row_reg, col_reg}<16'b0011100001110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100001110010) && ({row_reg, col_reg}<16'b0011100001110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011100001110100) && ({row_reg, col_reg}<16'b0011100001110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100001110110) && ({row_reg, col_reg}<16'b0011100001111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100001111001) && ({row_reg, col_reg}<16'b0011100001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100001111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100001111101) && ({row_reg, col_reg}<16'b0011100010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100010000011) && ({row_reg, col_reg}<16'b0011100010100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011100010100100) && ({row_reg, col_reg}<16'b0011100010100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100010100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100010100111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100010101000) && ({row_reg, col_reg}<16'b0011100010101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100010101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011100010101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011100010101110) && ({row_reg, col_reg}<16'b0011100010110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100010110001) && ({row_reg, col_reg}<16'b0011100010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011100010110011) && ({row_reg, col_reg}<16'b0011100010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100010110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100010110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011100010110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011100010111000) && ({row_reg, col_reg}<16'b0011100010111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100011000000) && ({row_reg, col_reg}<16'b0011100011000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011100011000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100011000011) && ({row_reg, col_reg}<16'b0011100011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100011001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100011001100) && ({row_reg, col_reg}<16'b0011100011001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011100011001110) && ({row_reg, col_reg}<16'b0011100011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100011011111) && ({row_reg, col_reg}<16'b0011100011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011100011100001) && ({row_reg, col_reg}<16'b0011100011100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100011100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100011100110) && ({row_reg, col_reg}<16'b0011100011101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011100011101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100011101001) && ({row_reg, col_reg}<16'b0011100011101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011100011101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100011101110) && ({row_reg, col_reg}<16'b0011100011110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011100011110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100011110001) && ({row_reg, col_reg}<16'b0011100011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011100011111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011100011111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100011111100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0011100011111101) && ({row_reg, col_reg}<16'b0011100100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011100100000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100100000001) && ({row_reg, col_reg}<16'b0011100100000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100100000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011100100000100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011100100000101)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0011100100000110) && ({row_reg, col_reg}<16'b0011100100001000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011100100001000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011100100001001)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=16'b0011100100001010) && ({row_reg, col_reg}<16'b0011100100001100)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011100100001100)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011100100001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011100100001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011100100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100100010000) && ({row_reg, col_reg}<16'b0011100100010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011100100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100100010011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011100100010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100100010101) && ({row_reg, col_reg}<16'b0011100100011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100100011001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011100100011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100100011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011100100011100) && ({row_reg, col_reg}<16'b0011100100011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011100100011111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011100100100000)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0011100100100001) && ({row_reg, col_reg}<16'b0011100100110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011100100110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011100100110001)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}>=16'b0011100100110010) && ({row_reg, col_reg}<16'b0011100100110100)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011100100110100)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011100100110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0011100100110110) && ({row_reg, col_reg}<16'b0011100100111000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011100100111000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0011100100111001) && ({row_reg, col_reg}<16'b0011100100111101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011100100111101)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0011100100111110) && ({row_reg, col_reg}<16'b0011100101000000)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}>=16'b0011100101000000) && ({row_reg, col_reg}<16'b0011100101000010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011100101000010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011100101000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011100101000100) && ({row_reg, col_reg}<16'b0011100101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100101000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011100101000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011100101001000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011100101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011100101001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011100101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011100101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100101001101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011100101001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011100101001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011100101010000) && ({row_reg, col_reg}<16'b0011100101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011100101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100101010101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0011100101010110) && ({row_reg, col_reg}<16'b0011100101011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100101011000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0011100101011001) && ({row_reg, col_reg}<16'b0011100101011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011100101011011) && ({row_reg, col_reg}<16'b0011100101011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011100101011101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011100101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100101011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100101100000) && ({row_reg, col_reg}<16'b0011100101100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011100101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100101100011) && ({row_reg, col_reg}<16'b0011100101100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100101100101) && ({row_reg, col_reg}<16'b0011100101100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011100101100111) && ({row_reg, col_reg}<16'b0011100101101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100101101001) && ({row_reg, col_reg}<16'b0011100101101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011100101101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011100101101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011100101101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011100101101110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0011100101101111) && ({row_reg, col_reg}<16'b0011100101110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011100101110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100101110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011100101110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011100101110100) && ({row_reg, col_reg}<16'b0011100101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100101110110) && ({row_reg, col_reg}<16'b0011100101111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100101111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100101111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100101111101) && ({row_reg, col_reg}<16'b0011100110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100110000011) && ({row_reg, col_reg}<16'b0011100110100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011100110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100110100101) && ({row_reg, col_reg}<16'b0011100110100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100110100111) && ({row_reg, col_reg}<16'b0011100110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100110101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100110101100) && ({row_reg, col_reg}<16'b0011100110101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011100110101110) && ({row_reg, col_reg}<16'b0011100110110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100110110000) && ({row_reg, col_reg}<16'b0011100110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011100110110011) && ({row_reg, col_reg}<16'b0011100110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100110110101) && ({row_reg, col_reg}<16'b0011100110110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100110110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100110111000) && ({row_reg, col_reg}<16'b0011100110111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100110111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011100110111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100110111100) && ({row_reg, col_reg}<16'b0011100110111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100110111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100111000000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==16'b0011100111000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011100111000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100111000011) && ({row_reg, col_reg}<16'b0011100111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100111001001) && ({row_reg, col_reg}<16'b0011100111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100111001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011100111001100) && ({row_reg, col_reg}<16'b0011100111010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011100111010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100111010001) && ({row_reg, col_reg}<16'b0011100111011101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011100111011101) && ({row_reg, col_reg}<16'b0011100111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100111011111) && ({row_reg, col_reg}<16'b0011100111100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011100111100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100111100010) && ({row_reg, col_reg}<16'b0011100111100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100111100100) && ({row_reg, col_reg}<16'b0011100111100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100111100110) && ({row_reg, col_reg}<16'b0011100111101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100111101000) && ({row_reg, col_reg}<16'b0011100111101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011100111101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100111101110) && ({row_reg, col_reg}<16'b0011100111110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011100111110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100111110001) && ({row_reg, col_reg}<16'b0011100111111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011100111111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011100111111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100111111100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0011100111111101) && ({row_reg, col_reg}<16'b0011101000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011101000000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101000000001) && ({row_reg, col_reg}<16'b0011101000000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101000000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011101000000100) && ({row_reg, col_reg}<16'b0011101000000110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011101000000110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0011101000000111) && ({row_reg, col_reg}<16'b0011101000001010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011101000001010)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0011101000001011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011101000001100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011101000001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011101000001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011101000001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011101000010000) && ({row_reg, col_reg}<16'b0011101000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011101000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101000010011) && ({row_reg, col_reg}<16'b0011101000010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101000010101) && ({row_reg, col_reg}<16'b0011101000011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011101000011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101000011001) && ({row_reg, col_reg}<16'b0011101000011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011101000011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101000011100) && ({row_reg, col_reg}<16'b0011101000011110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011101000011110) && ({row_reg, col_reg}<16'b0011101000100001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011101000100001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0011101000100010) && ({row_reg, col_reg}<16'b0011101000101111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011101000101111)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0011101000110000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011101000110001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0011101000110010) && ({row_reg, col_reg}<16'b0011101000110100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011101000110100)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0011101000110101) && ({row_reg, col_reg}<16'b0011101000111000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011101000111000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011101000111001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0011101000111010) && ({row_reg, col_reg}<16'b0011101000111101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011101000111101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0011101000111110) && ({row_reg, col_reg}<16'b0011101001000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011101001000000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011101001000001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011101001000010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011101001000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011101001000100) && ({row_reg, col_reg}<16'b0011101001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101001000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011101001000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011101001001000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011101001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011101001001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011101001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101001001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011101001001110) && ({row_reg, col_reg}<16'b0011101001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011101001010000) && ({row_reg, col_reg}<16'b0011101001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011101001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101001010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101001010110) && ({row_reg, col_reg}<16'b0011101001011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101001011000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0011101001011001) && ({row_reg, col_reg}<16'b0011101001011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011101001011011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011101001011100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011101001011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011101001011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011101001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101001100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011101001100001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011101001100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101001100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011101001100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011101001100101) && ({row_reg, col_reg}<16'b0011101001100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011101001100111) && ({row_reg, col_reg}<16'b0011101001101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101001101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011101001101011) && ({row_reg, col_reg}<16'b0011101001101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011101001101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011101001101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101001101111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0011101001110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011101001110001) && ({row_reg, col_reg}<16'b0011101001110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101001110011) && ({row_reg, col_reg}<16'b0011101001110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101001110110) && ({row_reg, col_reg}<16'b0011101010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101010000011) && ({row_reg, col_reg}<16'b0011101010100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011101010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101010100100) && ({row_reg, col_reg}<16'b0011101010100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011101010100111) && ({row_reg, col_reg}<16'b0011101010101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101010101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011101010101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011101010101110) && ({row_reg, col_reg}<16'b0011101010110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101010110000) && ({row_reg, col_reg}<16'b0011101010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011101010110011) && ({row_reg, col_reg}<16'b0011101010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011101010110101) && ({row_reg, col_reg}<16'b0011101010110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101010110111) && ({row_reg, col_reg}<16'b0011101010111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101010111001) && ({row_reg, col_reg}<16'b0011101010111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101010111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011101010111100) && ({row_reg, col_reg}<16'b0011101011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101011000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011101011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011101011000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101011000011) && ({row_reg, col_reg}<16'b0011101011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101011001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011101011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011101011001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011101011001100) && ({row_reg, col_reg}<16'b0011101011010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011101011010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101011010001) && ({row_reg, col_reg}<16'b0011101011011101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011101011011101) && ({row_reg, col_reg}<16'b0011101011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101011011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011101011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011101011100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101011100010) && ({row_reg, col_reg}<16'b0011101011100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101011100100) && ({row_reg, col_reg}<16'b0011101011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011101011100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101011101000) && ({row_reg, col_reg}<16'b0011101011101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011101011101100) && ({row_reg, col_reg}<16'b0011101011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101011101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011101011110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101011110001) && ({row_reg, col_reg}<16'b0011101011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011101011111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011101011111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101011111100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0011101011111101) && ({row_reg, col_reg}<16'b0011101100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011101100000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101100000001) && ({row_reg, col_reg}<16'b0011101100000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011101100000011) && ({row_reg, col_reg}<16'b0011101100000110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011101100000110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011101100000111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011101100001000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0011101100001001) && ({row_reg, col_reg}<16'b0011101100001011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0011101100001011) && ({row_reg, col_reg}<16'b0011101100001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011101100001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011101100001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011101100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011101100010000) && ({row_reg, col_reg}<16'b0011101100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011101100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101100010011) && ({row_reg, col_reg}<16'b0011101100010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101100010101) && ({row_reg, col_reg}<16'b0011101100011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011101100011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101100011001) && ({row_reg, col_reg}<16'b0011101100011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011101100011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101100011100) && ({row_reg, col_reg}<16'b0011101100011110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011101100011110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011101100011111) && ({row_reg, col_reg}<16'b0011101100100001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0011101100100001) && ({row_reg, col_reg}<16'b0011101100110001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011101100110001) && ({row_reg, col_reg}<16'b0011101100110011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011101100110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0011101100110100) && ({row_reg, col_reg}<16'b0011101100111010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011101100111010) && ({row_reg, col_reg}<16'b0011101100111101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011101100111101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011101100111110) && ({row_reg, col_reg}<16'b0011101101000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011101101000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011101101000001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011101101000010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011101101000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011101101000100) && ({row_reg, col_reg}<16'b0011101101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101101000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011101101000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011101101001000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011101101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011101101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101101001100) && ({row_reg, col_reg}<16'b0011101101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011101101010000) && ({row_reg, col_reg}<16'b0011101101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011101101010100) && ({row_reg, col_reg}<16'b0011101101011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011101101011000) && ({row_reg, col_reg}<16'b0011101101011011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011101101011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101101011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011101101011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011101101011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011101101011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101101100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101101100001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011101101100010) && ({row_reg, col_reg}<16'b0011101101100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101101100101) && ({row_reg, col_reg}<16'b0011101101100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011101101100111) && ({row_reg, col_reg}<16'b0011101101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101101101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011101101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011101101101100) && ({row_reg, col_reg}<16'b0011101101110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011101101110001) && ({row_reg, col_reg}<16'b0011101101110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101101110011) && ({row_reg, col_reg}<16'b0011101101110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101101110101) && ({row_reg, col_reg}<16'b0011101101111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101101111010) && ({row_reg, col_reg}<16'b0011101101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101101111111) && ({row_reg, col_reg}<16'b0011101110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101110000011) && ({row_reg, col_reg}<16'b0011101110100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011101110100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011101110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101110100101) && ({row_reg, col_reg}<16'b0011101110100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011101110100111) && ({row_reg, col_reg}<16'b0011101110101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101110101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101110101111) && ({row_reg, col_reg}<16'b0011101110110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011101110110001) && ({row_reg, col_reg}<16'b0011101110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011101110110011) && ({row_reg, col_reg}<16'b0011101110110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101110110111) && ({row_reg, col_reg}<16'b0011101110111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101110111001) && ({row_reg, col_reg}<16'b0011101110111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101110111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011101110111100) && ({row_reg, col_reg}<16'b0011101111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101111000000) && ({row_reg, col_reg}<16'b0011101111000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101111000011) && ({row_reg, col_reg}<16'b0011101111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101111001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011101111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101111001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011101111001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011101111001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011101111001101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0011101111001110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011101111001111) && ({row_reg, col_reg}<16'b0011101111011101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011101111011101) && ({row_reg, col_reg}<16'b0011101111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101111011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011101111100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011101111100001) && ({row_reg, col_reg}<16'b0011101111100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101111100100) && ({row_reg, col_reg}<16'b0011101111100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011101111100111) && ({row_reg, col_reg}<16'b0011101111101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101111101001) && ({row_reg, col_reg}<16'b0011101111101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011101111101101) && ({row_reg, col_reg}<16'b0011101111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101111110001) && ({row_reg, col_reg}<16'b0011101111111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011101111111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011101111111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101111111100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0011101111111101) && ({row_reg, col_reg}<16'b0011110000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011110000000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110000000001) && ({row_reg, col_reg}<16'b0011110000000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110000000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011110000000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011110000000101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011110000000110) && ({row_reg, col_reg}<16'b0011110000001000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011110000001000) && ({row_reg, col_reg}<16'b0011110000001010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011110000001010)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}>=16'b0011110000001011) && ({row_reg, col_reg}<16'b0011110000001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011110000001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011110000001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011110000001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110000010000) && ({row_reg, col_reg}<16'b0011110000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110000010010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011110000010011) && ({row_reg, col_reg}<16'b0011110000010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110000010101) && ({row_reg, col_reg}<16'b0011110000011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011110000011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110000011001) && ({row_reg, col_reg}<16'b0011110000011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011110000011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110000011100) && ({row_reg, col_reg}<16'b0011110000011110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011110000011110) && ({row_reg, col_reg}<16'b0011110000100000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011110000100000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0011110000100001) && ({row_reg, col_reg}<16'b0011110000110101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011110000110101)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0011110000110110) && ({row_reg, col_reg}<16'b0011110000111000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011110000111000) && ({row_reg, col_reg}<16'b0011110000111011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011110000111011)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0011110000111100) && ({row_reg, col_reg}<16'b0011110000111110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011110000111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011110000111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011110001000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011110001000001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011110001000010)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0011110001000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011110001000100) && ({row_reg, col_reg}<16'b0011110001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110001000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011110001000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011110001001000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011110001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011110001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110001001100) && ({row_reg, col_reg}<16'b0011110001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011110001010000) && ({row_reg, col_reg}<16'b0011110001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011110001010100) && ({row_reg, col_reg}<16'b0011110001011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110001011000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011110001011001) && ({row_reg, col_reg}<16'b0011110001011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110001011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011110001011110) && ({row_reg, col_reg}<16'b0011110001100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011110001100000) && ({row_reg, col_reg}<16'b0011110001100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110001100101) && ({row_reg, col_reg}<16'b0011110001101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011110001101010) && ({row_reg, col_reg}<16'b0011110001101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110001101100) && ({row_reg, col_reg}<16'b0011110001110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011110001110001) && ({row_reg, col_reg}<16'b0011110001111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110001111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011110001111011) && ({row_reg, col_reg}<16'b0011110010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110010000000) && ({row_reg, col_reg}<16'b0011110010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110010000011) && ({row_reg, col_reg}<16'b0011110010100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011110010100100) && ({row_reg, col_reg}<16'b0011110010100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110010100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011110010101000) && ({row_reg, col_reg}<16'b0011110010101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110010101010) && ({row_reg, col_reg}<16'b0011110010101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110010101100) && ({row_reg, col_reg}<16'b0011110010101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110010101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110010101111) && ({row_reg, col_reg}<16'b0011110010110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110010110001) && ({row_reg, col_reg}<16'b0011110010110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110010110100) && ({row_reg, col_reg}<16'b0011110010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110010110110) && ({row_reg, col_reg}<16'b0011110010111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110010111001) && ({row_reg, col_reg}<16'b0011110011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110011000000) && ({row_reg, col_reg}<16'b0011110011000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110011000011) && ({row_reg, col_reg}<16'b0011110011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110011001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011110011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110011001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011110011001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011110011001101) && ({row_reg, col_reg}<16'b0011110011001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011110011001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011110011010000) && ({row_reg, col_reg}<16'b0011110011010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110011010010) && ({row_reg, col_reg}<16'b0011110011011101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011110011011101) && ({row_reg, col_reg}<16'b0011110011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110011011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011110011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011110011100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110011100010) && ({row_reg, col_reg}<16'b0011110011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110011100111) && ({row_reg, col_reg}<16'b0011110011101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110011101010) && ({row_reg, col_reg}<16'b0011110011101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011110011101101) && ({row_reg, col_reg}<16'b0011110011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110011101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110011110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110011110001) && ({row_reg, col_reg}<16'b0011110011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011110011111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011110011111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110011111100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0011110011111101) && ({row_reg, col_reg}<16'b0011110100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011110100000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110100000001) && ({row_reg, col_reg}<16'b0011110100000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011110100000011) && ({row_reg, col_reg}<16'b0011110100000101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011110100000101)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0011110100000110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011110100000111) && ({row_reg, col_reg}<16'b0011110100001010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011110100001010)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}>=16'b0011110100001011) && ({row_reg, col_reg}<16'b0011110100001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011110100001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011110100001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011110100001111) && ({row_reg, col_reg}<16'b0011110100010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110100010101) && ({row_reg, col_reg}<16'b0011110100011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011110100011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110100011001) && ({row_reg, col_reg}<16'b0011110100011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011110100011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110100011100) && ({row_reg, col_reg}<16'b0011110100011110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011110100011110) && ({row_reg, col_reg}<16'b0011110100100000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011110100100000) && ({row_reg, col_reg}<16'b0011110100110001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0011110100110001) && ({row_reg, col_reg}<16'b0011110100110011)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0011110100110011)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0011110100110100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011110100110101)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0011110100110110) && ({row_reg, col_reg}<16'b0011110100111101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011110100111101) && ({row_reg, col_reg}<16'b0011110101000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011110101000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011110101000001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0011110101000010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011110101000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011110101000100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011110101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110101000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011110101000111) && ({row_reg, col_reg}<16'b0011110101001001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011110101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011110101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110101001100) && ({row_reg, col_reg}<16'b0011110101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011110101010000) && ({row_reg, col_reg}<16'b0011110101010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011110101010010)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0011110101010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011110101010100) && ({row_reg, col_reg}<16'b0011110101010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110101010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110101010111) && ({row_reg, col_reg}<16'b0011110101011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110101011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011110101100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011110101100001) && ({row_reg, col_reg}<16'b0011110101100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011110101100011) && ({row_reg, col_reg}<16'b0011110101100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110101100101) && ({row_reg, col_reg}<16'b0011110101100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011110101100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011110101101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011110101101001)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b0011110101101010) && ({row_reg, col_reg}<16'b0011110101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110101101100) && ({row_reg, col_reg}<16'b0011110101101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011110101101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011110101110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110101110001) && ({row_reg, col_reg}<16'b0011110101110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110101110011) && ({row_reg, col_reg}<16'b0011110101110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110101110101) && ({row_reg, col_reg}<16'b0011110101111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110101111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110101111010) && ({row_reg, col_reg}<16'b0011110101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011110101111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110101111101) && ({row_reg, col_reg}<16'b0011110101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110110000000) && ({row_reg, col_reg}<16'b0011110110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110110000011) && ({row_reg, col_reg}<16'b0011110110100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011110110100100) && ({row_reg, col_reg}<16'b0011110110100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110110100110) && ({row_reg, col_reg}<16'b0011110110101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011110110101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110110101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110110101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011110110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110110101100) && ({row_reg, col_reg}<16'b0011110110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110110110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110110110001) && ({row_reg, col_reg}<16'b0011110110110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110110110011) && ({row_reg, col_reg}<16'b0011110110110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110110110101) && ({row_reg, col_reg}<16'b0011110110110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011110110110111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=16'b0011110110111000) && ({row_reg, col_reg}<16'b0011110111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110111000000) && ({row_reg, col_reg}<16'b0011110111000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011110111000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110111000011) && ({row_reg, col_reg}<16'b0011110111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110111001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011110111001001) && ({row_reg, col_reg}<16'b0011110111001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110111001011) && ({row_reg, col_reg}<16'b0011110111001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011110111001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011110111001110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011110111001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011110111010000) && ({row_reg, col_reg}<16'b0011110111010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110111010010) && ({row_reg, col_reg}<16'b0011110111010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011110111010100) && ({row_reg, col_reg}<16'b0011110111011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110111011000) && ({row_reg, col_reg}<16'b0011110111011101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011110111011101) && ({row_reg, col_reg}<16'b0011110111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110111011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011110111100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011110111100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011110111100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110111100011) && ({row_reg, col_reg}<16'b0011110111100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110111100111) && ({row_reg, col_reg}<16'b0011110111101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110111101001) && ({row_reg, col_reg}<16'b0011110111101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011110111101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110111101110) && ({row_reg, col_reg}<16'b0011110111110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110111110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110111110001) && ({row_reg, col_reg}<16'b0011110111111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011110111111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011110111111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110111111100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0011110111111101) && ({row_reg, col_reg}<16'b0011111000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111000000000) && ({row_reg, col_reg}<16'b0011111000000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011111000000011) && ({row_reg, col_reg}<16'b0011111000000110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111000000110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011111000000111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0011111000001000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011111000001001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011111000001010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011111000001011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011111000001100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111000001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011111000001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111000001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011111000010000) && ({row_reg, col_reg}<16'b0011111000010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111000010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011111000010011) && ({row_reg, col_reg}<16'b0011111000010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011111000010101) && ({row_reg, col_reg}<16'b0011111000011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111000011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011111000011001) && ({row_reg, col_reg}<16'b0011111000011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011111000011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011111000011100) && ({row_reg, col_reg}<16'b0011111000011110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011111000011110) && ({row_reg, col_reg}<16'b0011111000100000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011111000100000)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0011111000100001) && ({row_reg, col_reg}<16'b0011111000110111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011111000110111) && ({row_reg, col_reg}<16'b0011111000111001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0011111000111001) && ({row_reg, col_reg}<16'b0011111000111100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011111000111100) && ({row_reg, col_reg}<16'b0011111000111110)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0011111000111110) && ({row_reg, col_reg}<16'b0011111001000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011111001000000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011111001000001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011111001000010)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0011111001000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011111001000100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011111001000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011111001000110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0011111001000111) && ({row_reg, col_reg}<16'b0011111001001001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011111001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011111001001010) && ({row_reg, col_reg}<16'b0011111001001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111001001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011111001001110) && ({row_reg, col_reg}<16'b0011111001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011111001010000) && ({row_reg, col_reg}<16'b0011111001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011111001010100) && ({row_reg, col_reg}<16'b0011111001010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111001010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011111001010111) && ({row_reg, col_reg}<16'b0011111001011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011111001011110) && ({row_reg, col_reg}<16'b0011111001100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111001100000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011111001100001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111001100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111001100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011111001100101) && ({row_reg, col_reg}<16'b0011111001100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011111001100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111001101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011111001101001)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}>=16'b0011111001101010) && ({row_reg, col_reg}<16'b0011111001101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011111001101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011111001101101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0011111001101110) && ({row_reg, col_reg}<16'b0011111001110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111001110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111001110001) && ({row_reg, col_reg}<16'b0011111001110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111001110101) && ({row_reg, col_reg}<16'b0011111001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011111001111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011111001111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111001111101) && ({row_reg, col_reg}<16'b0011111001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111010000000) && ({row_reg, col_reg}<16'b0011111010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111010000011) && ({row_reg, col_reg}<16'b0011111010100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011111010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111010100100) && ({row_reg, col_reg}<16'b0011111010100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111010100110) && ({row_reg, col_reg}<16'b0011111010101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111010101000) && ({row_reg, col_reg}<16'b0011111010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111010101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111010101011) && ({row_reg, col_reg}<16'b0011111010101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111010101111) && ({row_reg, col_reg}<16'b0011111010110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111010110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111010110010) && ({row_reg, col_reg}<16'b0011111010110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111010110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011111010110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111010110110) && ({row_reg, col_reg}<16'b0011111010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111010111000) && ({row_reg, col_reg}<16'b0011111010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111010111110) && ({row_reg, col_reg}<16'b0011111011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111011000000) && ({row_reg, col_reg}<16'b0011111011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111011000011) && ({row_reg, col_reg}<16'b0011111011000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111011000101) && ({row_reg, col_reg}<16'b0011111011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111011001000) && ({row_reg, col_reg}<16'b0011111011010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011111011010100) && ({row_reg, col_reg}<16'b0011111011011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111011011001) && ({row_reg, col_reg}<16'b0011111011011101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011111011011101) && ({row_reg, col_reg}<16'b0011111011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111011011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011111011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011111011100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111011100010) && ({row_reg, col_reg}<16'b0011111011100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111011100100) && ({row_reg, col_reg}<16'b0011111011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111011100111) && ({row_reg, col_reg}<16'b0011111011101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111011101001) && ({row_reg, col_reg}<16'b0011111011101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011111011101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111011101110) && ({row_reg, col_reg}<16'b0011111011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011111011110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111011110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111011110010) && ({row_reg, col_reg}<16'b0011111011111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011111011111011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0011111011111100) && ({row_reg, col_reg}<16'b0011111100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111100000000) && ({row_reg, col_reg}<16'b0011111100000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111100000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111100000100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0011111100000101) && ({row_reg, col_reg}<16'b0011111100000111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011111100000111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0011111100001000) && ({row_reg, col_reg}<16'b0011111100001011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0011111100001011) && ({row_reg, col_reg}<16'b0011111100001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011111100001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111100001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011111100001111) && ({row_reg, col_reg}<16'b0011111100010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011111100010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111100010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011111100010011) && ({row_reg, col_reg}<16'b0011111100010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011111100010101) && ({row_reg, col_reg}<16'b0011111100011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111100011000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011111100011001) && ({row_reg, col_reg}<16'b0011111100011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111100011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011111100011100) && ({row_reg, col_reg}<16'b0011111100011110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111100011110)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0011111100011111) && ({row_reg, col_reg}<16'b0011111100110101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011111100110101)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0011111100110110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011111100110111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0011111100111000) && ({row_reg, col_reg}<16'b0011111100111100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011111100111100) && ({row_reg, col_reg}<16'b0011111100111110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011111100111110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011111100111111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0011111101000000)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011111101000001)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011111101000010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011111101000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011111101000100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011111101000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011111101000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011111101000111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011111101001000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011111101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011111101001010) && ({row_reg, col_reg}<16'b0011111101001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111101001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011111101001110) && ({row_reg, col_reg}<16'b0011111101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011111101010000) && ({row_reg, col_reg}<16'b0011111101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011111101010100) && ({row_reg, col_reg}<16'b0011111101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011111101011110) && ({row_reg, col_reg}<16'b0011111101100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011111101100000) && ({row_reg, col_reg}<16'b0011111101100010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111101100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111101100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011111101100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111101100101) && ({row_reg, col_reg}<16'b0011111101100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011111101100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011111101101000) && ({row_reg, col_reg}<16'b0011111101101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011111101101010)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==16'b0011111101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011111101101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011111101101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111101101110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011111101101111) && ({row_reg, col_reg}<16'b0011111101110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011111101110001) && ({row_reg, col_reg}<16'b0011111101110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011111101110011) && ({row_reg, col_reg}<16'b0011111101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011111101111011)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=16'b0011111101111100) && ({row_reg, col_reg}<16'b0011111110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111110000000) && ({row_reg, col_reg}<16'b0011111110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111110000010) && ({row_reg, col_reg}<16'b0011111110100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011111110100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011111110100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111110100100) && ({row_reg, col_reg}<16'b0011111110100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111110100110) && ({row_reg, col_reg}<16'b0011111110101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011111110101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011111110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111110101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111110101011) && ({row_reg, col_reg}<16'b0011111110101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111110101110) && ({row_reg, col_reg}<16'b0011111110110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111110110110) && ({row_reg, col_reg}<16'b0011111110111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111110111001) && ({row_reg, col_reg}<16'b0011111110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111110111101) && ({row_reg, col_reg}<16'b0011111111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011111111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111111000001) && ({row_reg, col_reg}<16'b0011111111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111111000011) && ({row_reg, col_reg}<16'b0011111111000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111111000101) && ({row_reg, col_reg}<16'b0011111111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111111000111) && ({row_reg, col_reg}<16'b0011111111010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011111111010100) && ({row_reg, col_reg}<16'b0011111111011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111111011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011111111011101) && ({row_reg, col_reg}<16'b0011111111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111111011111) && ({row_reg, col_reg}<16'b0011111111100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011111111100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011111111100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111111100011) && ({row_reg, col_reg}<16'b0011111111100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111111100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111111100111) && ({row_reg, col_reg}<16'b0011111111101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111111101001) && ({row_reg, col_reg}<16'b0011111111101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011111111101101) && ({row_reg, col_reg}<16'b0011111111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111111101111) && ({row_reg, col_reg}<16'b0011111111110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011111111110001)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0011111111110010) && ({row_reg, col_reg}<16'b0100000000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000000000000) && ({row_reg, col_reg}<16'b0100000000000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000000000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000000000100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100000000000101)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100000000000110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100000000000111) && ({row_reg, col_reg}<16'b0100000000001010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100000000001010)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100000000001011) && ({row_reg, col_reg}<16'b0100000000001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100000000001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000000001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100000000001111) && ({row_reg, col_reg}<16'b0100000000010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100000000010101) && ({row_reg, col_reg}<16'b0100000000011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000000011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100000000011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000000011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100000000011100) && ({row_reg, col_reg}<16'b0100000000011110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000000011110)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0100000000011111) && ({row_reg, col_reg}<16'b0100000000110011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100000000110011) && ({row_reg, col_reg}<16'b0100000000110101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100000000110101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100000000110110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100000000110111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100000000111000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100000000111001)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0100000000111010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000000111011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100000000111100)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100000000111101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100000000111110) && ({row_reg, col_reg}<16'b0100000001000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100000001000000)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0100000001000001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0100000001000010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0100000001000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100000001000100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100000001000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100000001000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100000001000111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100000001001000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100000001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100000001001010) && ({row_reg, col_reg}<16'b0100000001001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000001001101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0100000001001110) && ({row_reg, col_reg}<16'b0100000001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000001010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100000001010001) && ({row_reg, col_reg}<16'b0100000001010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000001010011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0100000001010100) && ({row_reg, col_reg}<16'b0100000001010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100000001010111) && ({row_reg, col_reg}<16'b0100000001011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100000001011110) && ({row_reg, col_reg}<16'b0100000001100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100000001100000) && ({row_reg, col_reg}<16'b0100000001100010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000001100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100000001100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100000001100101) && ({row_reg, col_reg}<16'b0100000001100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100000001100111) && ({row_reg, col_reg}<16'b0100000001101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100000001101001) && ({row_reg, col_reg}<16'b0100000001101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100000001101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000001101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100000001101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100000001101110) && ({row_reg, col_reg}<16'b0100000001110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000001110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100000001110001) && ({row_reg, col_reg}<16'b0100000001110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100000001110011) && ({row_reg, col_reg}<16'b0100000001111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100000001111001) && ({row_reg, col_reg}<16'b0100000001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000001111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000001111101) && ({row_reg, col_reg}<16'b0100000010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000010000000) && ({row_reg, col_reg}<16'b0100000010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000010000011) && ({row_reg, col_reg}<16'b0100000010100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100000010100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100000010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000010100100) && ({row_reg, col_reg}<16'b0100000010100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100000010100110) && ({row_reg, col_reg}<16'b0100000010101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100000010101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100000010101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000010101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000010101011) && ({row_reg, col_reg}<16'b0100000010101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100000010101101) && ({row_reg, col_reg}<16'b0100000010110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000010110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000010110010) && ({row_reg, col_reg}<16'b0100000010110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000010110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100000010110101) && ({row_reg, col_reg}<16'b0100000010110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000010110111) && ({row_reg, col_reg}<16'b0100000010111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000010111001) && ({row_reg, col_reg}<16'b0100000010111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000010111101) && ({row_reg, col_reg}<16'b0100000011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100000011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000011000001) && ({row_reg, col_reg}<16'b0100000011000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000011000101) && ({row_reg, col_reg}<16'b0100000011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000011001000) && ({row_reg, col_reg}<16'b0100000011001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100000011001100) && ({row_reg, col_reg}<16'b0100000011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000011001110) && ({row_reg, col_reg}<16'b0100000011010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100000011010011) && ({row_reg, col_reg}<16'b0100000011011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000011011100) && ({row_reg, col_reg}<16'b0100000011011110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100000011011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000011011111) && ({row_reg, col_reg}<16'b0100000011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100000011100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000011100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100000011100011) && ({row_reg, col_reg}<16'b0100000011100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000011100110) && ({row_reg, col_reg}<16'b0100000011101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100000011101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000011101001) && ({row_reg, col_reg}<16'b0100000011101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100000011101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100000011110000)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0100000011110001) && ({row_reg, col_reg}<16'b0100000100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000100000000) && ({row_reg, col_reg}<16'b0100000100000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000100000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100000100000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0100000100000101) && ({row_reg, col_reg}<16'b0100000100000111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100000100000111) && ({row_reg, col_reg}<16'b0100000100001001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100000100001001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0100000100001010) && ({row_reg, col_reg}<16'b0100000100001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100000100001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000100001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000100001111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100000100010000) && ({row_reg, col_reg}<16'b0100000100010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000100010011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100000100010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100000100010101) && ({row_reg, col_reg}<16'b0100000100011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000100011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000100011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100000100011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100000100011100) && ({row_reg, col_reg}<16'b0100000100011110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000100011110)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0100000100011111) && ({row_reg, col_reg}<16'b0100000100110100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000100110100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100000100110101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100000100110110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100000100110111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100000100111000) && ({row_reg, col_reg}<16'b0100000100111100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100000100111100) && ({row_reg, col_reg}<16'b0100000100111110)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100000100111110) && ({row_reg, col_reg}<16'b0100000101000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100000101000000)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0100000101000001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0100000101000010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0100000101000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100000101000100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100000101000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100000101000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100000101000111)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0100000101001000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100000101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100000101001010) && ({row_reg, col_reg}<16'b0100000101001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100000101001101) && ({row_reg, col_reg}<16'b0100000101001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100000101001111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000101010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100000101010001) && ({row_reg, col_reg}<16'b0100000101010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100000101010011) && ({row_reg, col_reg}<16'b0100000101010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100000101010111) && ({row_reg, col_reg}<16'b0100000101011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100000101011100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0100000101011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100000101011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0100000101011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100000101100000) && ({row_reg, col_reg}<16'b0100000101100010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100000101100011) && ({row_reg, col_reg}<16'b0100000101100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100000101100101) && ({row_reg, col_reg}<16'b0100000101101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100000101101000) && ({row_reg, col_reg}<16'b0100000101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000101101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100000101101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100000101101100) && ({row_reg, col_reg}<16'b0100000101101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100000101101110) && ({row_reg, col_reg}<16'b0100000101110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100000101110001) && ({row_reg, col_reg}<16'b0100000101110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000101110011) && ({row_reg, col_reg}<16'b0100000101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100000101110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000101110111) && ({row_reg, col_reg}<16'b0100000101111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100000101111001) && ({row_reg, col_reg}<16'b0100000101111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000101111100) && ({row_reg, col_reg}<16'b0100000110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000110000000) && ({row_reg, col_reg}<16'b0100000110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000110000011) && ({row_reg, col_reg}<16'b0100000110100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100000110100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100000110100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000110100100) && ({row_reg, col_reg}<16'b0100000110100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100000110100110) && ({row_reg, col_reg}<16'b0100000110101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000110101000) && ({row_reg, col_reg}<16'b0100000110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000110101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100000110101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000110101100) && ({row_reg, col_reg}<16'b0100000110110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000110110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000110110010) && ({row_reg, col_reg}<16'b0100000110110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000110110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100000110110101) && ({row_reg, col_reg}<16'b0100000110110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000110110111) && ({row_reg, col_reg}<16'b0100000110111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000110111001) && ({row_reg, col_reg}<16'b0100000110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000110111101) && ({row_reg, col_reg}<16'b0100000111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100000111000000) && ({row_reg, col_reg}<16'b0100000111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000111000011) && ({row_reg, col_reg}<16'b0100000111000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000111000101) && ({row_reg, col_reg}<16'b0100000111001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000111001010) && ({row_reg, col_reg}<16'b0100000111001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100000111001100) && ({row_reg, col_reg}<16'b0100000111001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000111001111) && ({row_reg, col_reg}<16'b0100000111010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100000111010010) && ({row_reg, col_reg}<16'b0100000111011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000111011010) && ({row_reg, col_reg}<16'b0100000111011101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100000111011101) && ({row_reg, col_reg}<16'b0100000111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000111011111) && ({row_reg, col_reg}<16'b0100000111100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100000111100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000111100010) && ({row_reg, col_reg}<16'b0100000111100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000111100100) && ({row_reg, col_reg}<16'b0100000111100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100000111100111) && ({row_reg, col_reg}<16'b0100000111101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000111101001) && ({row_reg, col_reg}<16'b0100000111101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100000111101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100000111110000)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0100000111110001) && ({row_reg, col_reg}<16'b0100001000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100001000000000) && ({row_reg, col_reg}<16'b0100001000000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001000000011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100001000000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100001000000101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100001000000110)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}>=16'b0100001000000111) && ({row_reg, col_reg}<16'b0100001000001001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100001000001001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100001000001010) && ({row_reg, col_reg}<16'b0100001000001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100001000001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100001000001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100001000001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001000010000) && ({row_reg, col_reg}<16'b0100001000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100001000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001000010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100001000010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001000010101) && ({row_reg, col_reg}<16'b0100001000011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100001000011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100001000011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100001000011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001000011100) && ({row_reg, col_reg}<16'b0100001000011110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100001000011110) && ({row_reg, col_reg}<16'b0100001000100000)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0100001000100000) && ({row_reg, col_reg}<16'b0100001000100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100001000100110) && ({row_reg, col_reg}<16'b0100001000101010)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0100001000101010) && ({row_reg, col_reg}<16'b0100001000101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100001000101101) && ({row_reg, col_reg}<16'b0100001000110000)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0100001000110000)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0100001000110001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100001000110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100001000110011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100001000110100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100001000110101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100001000110110) && ({row_reg, col_reg}<16'b0100001000111001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100001000111001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100001000111010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100001000111011)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100001000111100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100001000111101)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100001000111110) && ({row_reg, col_reg}<16'b0100001001000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100001001000000)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0100001001000001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0100001001000010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0100001001000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001001000100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100001001000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100001001000110) && ({row_reg, col_reg}<16'b0100001001001001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100001001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100001001001100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100001001001101) && ({row_reg, col_reg}<16'b0100001001010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100001001010000) && ({row_reg, col_reg}<16'b0100001001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100001001010100) && ({row_reg, col_reg}<16'b0100001001011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001001011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100001001011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001001011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0100001001011111) && ({row_reg, col_reg}<16'b0100001001100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001001100001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100001001100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001001100011) && ({row_reg, col_reg}<16'b0100001001100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100001001100101) && ({row_reg, col_reg}<16'b0100001001101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100001001101000) && ({row_reg, col_reg}<16'b0100001001101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001001101010) && ({row_reg, col_reg}<16'b0100001001101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100001001101100) && ({row_reg, col_reg}<16'b0100001001101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100001001101110) && ({row_reg, col_reg}<16'b0100001001110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100001001110000) && ({row_reg, col_reg}<16'b0100001001110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001001110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001001110011) && ({row_reg, col_reg}<16'b0100001001110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100001001110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001001110110) && ({row_reg, col_reg}<16'b0100001001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001001111111) && ({row_reg, col_reg}<16'b0100001010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100001010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001010000011) && ({row_reg, col_reg}<16'b0100001010100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100001010100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001010100011) && ({row_reg, col_reg}<16'b0100001010100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001010100111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001010101000) && ({row_reg, col_reg}<16'b0100001010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001010101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100001010101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100001010101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001010101101) && ({row_reg, col_reg}<16'b0100001010110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001010110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001010110010) && ({row_reg, col_reg}<16'b0100001010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001010110110) && ({row_reg, col_reg}<16'b0100001010111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001010111001) && ({row_reg, col_reg}<16'b0100001010111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001010111101) && ({row_reg, col_reg}<16'b0100001011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001011000000) && ({row_reg, col_reg}<16'b0100001011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100001011000011) && ({row_reg, col_reg}<16'b0100001011000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001011000101) && ({row_reg, col_reg}<16'b0100001011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001011001010) && ({row_reg, col_reg}<16'b0100001011010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100001011010010) && ({row_reg, col_reg}<16'b0100001011011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001011011001) && ({row_reg, col_reg}<16'b0100001011011101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100001011011101) && ({row_reg, col_reg}<16'b0100001011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001011011111) && ({row_reg, col_reg}<16'b0100001011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100001011100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001011100010) && ({row_reg, col_reg}<16'b0100001011100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001011100100) && ({row_reg, col_reg}<16'b0100001011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001011100111) && ({row_reg, col_reg}<16'b0100001011101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001011101010) && ({row_reg, col_reg}<16'b0100001011101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100001011101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001011101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100001011101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100001011110000)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0100001011110001) && ({row_reg, col_reg}<16'b0100001100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100001100000000) && ({row_reg, col_reg}<16'b0100001100000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001100000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001100000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100001100000101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100001100000110)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}>=16'b0100001100000111) && ({row_reg, col_reg}<16'b0100001100001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100001100001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100001100001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100001100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001100010000) && ({row_reg, col_reg}<16'b0100001100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100001100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001100010011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100001100010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001100010101) && ({row_reg, col_reg}<16'b0100001100011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100001100011001) && ({row_reg, col_reg}<16'b0100001100011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100001100011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100001100011100) && ({row_reg, col_reg}<16'b0100001100011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100001100011111)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0100001100100000) && ({row_reg, col_reg}<16'b0100001100100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100001100100110) && ({row_reg, col_reg}<16'b0100001100101000)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0100001100101000)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0100001100101001) && ({row_reg, col_reg}<16'b0100001100101101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100001100101101) && ({row_reg, col_reg}<16'b0100001100110000)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0100001100110000)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0100001100110001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100001100110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100001100110011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100001100110100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100001100110101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100001100110110) && ({row_reg, col_reg}<16'b0100001100111001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100001100111001) && ({row_reg, col_reg}<16'b0100001100111011)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100001100111011) && ({row_reg, col_reg}<16'b0100001100111101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100001100111101)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100001100111110) && ({row_reg, col_reg}<16'b0100001101000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100001101000000)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0100001101000001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0100001101000010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0100001101000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100001101000100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0100001101000101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0100001101000110) && ({row_reg, col_reg}<16'b0100001101001000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100001101001000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100001101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100001101001010) && ({row_reg, col_reg}<16'b0100001101001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100001101001100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100001101001101) && ({row_reg, col_reg}<16'b0100001101010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100001101010000) && ({row_reg, col_reg}<16'b0100001101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100001101010100) && ({row_reg, col_reg}<16'b0100001101011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001101011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100001101011110) && ({row_reg, col_reg}<16'b0100001101100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001101100011) && ({row_reg, col_reg}<16'b0100001101100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100001101100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100001101100110)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==16'b0100001101100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100001101101000) && ({row_reg, col_reg}<16'b0100001101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100001101101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100001101101011)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}>=16'b0100001101101100) && ({row_reg, col_reg}<16'b0100001101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001101101111) && ({row_reg, col_reg}<16'b0100001101110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001101110010) && ({row_reg, col_reg}<16'b0100001101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001101110110) && ({row_reg, col_reg}<16'b0100001101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001101111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001101111001) && ({row_reg, col_reg}<16'b0100001110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001110000011) && ({row_reg, col_reg}<16'b0100001110100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100001110100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001110100011) && ({row_reg, col_reg}<16'b0100001110100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001110100101) && ({row_reg, col_reg}<16'b0100001110101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001110101000) && ({row_reg, col_reg}<16'b0100001110101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001110101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001110101101) && ({row_reg, col_reg}<16'b0100001110110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001110110010) && ({row_reg, col_reg}<16'b0100001110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100001110110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100001110110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001110111000) && ({row_reg, col_reg}<16'b0100001110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001110111110) && ({row_reg, col_reg}<16'b0100001111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001111000000) && ({row_reg, col_reg}<16'b0100001111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100001111000011) && ({row_reg, col_reg}<16'b0100001111000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001111000101) && ({row_reg, col_reg}<16'b0100001111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001111001001) && ({row_reg, col_reg}<16'b0100001111010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100001111010011) && ({row_reg, col_reg}<16'b0100001111011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001111011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100001111011101) && ({row_reg, col_reg}<16'b0100001111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001111011111) && ({row_reg, col_reg}<16'b0100001111100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100001111100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001111100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001111100100) && ({row_reg, col_reg}<16'b0100001111100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001111100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001111100111) && ({row_reg, col_reg}<16'b0100001111101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001111101010) && ({row_reg, col_reg}<16'b0100001111101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100001111101101) && ({row_reg, col_reg}<16'b0100001111110001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0100001111110001) && ({row_reg, col_reg}<16'b0100010000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010000000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010000000001) && ({row_reg, col_reg}<16'b0100010000000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010000000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100010000000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100010000000101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100010000000110)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0100010000000111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100010000001000)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100010000001001) && ({row_reg, col_reg}<16'b0100010000001011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100010000001011) && ({row_reg, col_reg}<16'b0100010000001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100010000001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100010000001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100010000001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010000010000) && ({row_reg, col_reg}<16'b0100010000010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010000010011) && ({row_reg, col_reg}<16'b0100010000010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010000010101) && ({row_reg, col_reg}<16'b0100010000011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100010000011001) && ({row_reg, col_reg}<16'b0100010000011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100010000011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100010000011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100010000011110) && ({row_reg, col_reg}<16'b0100010000100001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100010000100001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100010000100010) && ({row_reg, col_reg}<16'b0100010000100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010000100100) && ({row_reg, col_reg}<16'b0100010000101010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100010000101010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100010000101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100010000101100) && ({row_reg, col_reg}<16'b0100010000110001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100010000110001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100010000110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100010000110011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100010000110100)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100010000110101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100010000110110)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100010000110111) && ({row_reg, col_reg}<16'b0100010000111001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100010000111001)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0100010000111010) && ({row_reg, col_reg}<16'b0100010000111101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100010000111101)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100010000111110) && ({row_reg, col_reg}<16'b0100010001000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100010001000000)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0100010001000001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0100010001000010)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}>=16'b0100010001000011) && ({row_reg, col_reg}<16'b0100010001000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100010001000101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0100010001000110) && ({row_reg, col_reg}<16'b0100010001001000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100010001001000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100010001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100010001001010) && ({row_reg, col_reg}<16'b0100010001001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010001001100) && ({row_reg, col_reg}<16'b0100010001001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100010001001111) && ({row_reg, col_reg}<16'b0100010001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100010001010100) && ({row_reg, col_reg}<16'b0100010001011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100010001011010) && ({row_reg, col_reg}<16'b0100010001011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100010001011101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0100010001011110) && ({row_reg, col_reg}<16'b0100010001100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100010001100011) && ({row_reg, col_reg}<16'b0100010001100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010001100101) && ({row_reg, col_reg}<16'b0100010001100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100010001100111) && ({row_reg, col_reg}<16'b0100010001101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010001101100) && ({row_reg, col_reg}<16'b0100010001101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010001101111) && ({row_reg, col_reg}<16'b0100010001110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010001110011) && ({row_reg, col_reg}<16'b0100010001110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100010001110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010001110111) && ({row_reg, col_reg}<16'b0100010001111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010001111001) && ({row_reg, col_reg}<16'b0100010001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010001111101) && ({row_reg, col_reg}<16'b0100010001111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010001111111) && ({row_reg, col_reg}<16'b0100010010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010010000011) && ({row_reg, col_reg}<16'b0100010010100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010010100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010010100011) && ({row_reg, col_reg}<16'b0100010010100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010010100101) && ({row_reg, col_reg}<16'b0100010010100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010010100111) && ({row_reg, col_reg}<16'b0100010010101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010010101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010010101101) && ({row_reg, col_reg}<16'b0100010010110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010010110001) && ({row_reg, col_reg}<16'b0100010010110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010010110100) && ({row_reg, col_reg}<16'b0100010010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010010110110) && ({row_reg, col_reg}<16'b0100010010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100010010111000) && ({row_reg, col_reg}<16'b0100010010111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010010111110) && ({row_reg, col_reg}<16'b0100010011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010011000000) && ({row_reg, col_reg}<16'b0100010011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100010011000011) && ({row_reg, col_reg}<16'b0100010011000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010011000101) && ({row_reg, col_reg}<16'b0100010011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010011001001) && ({row_reg, col_reg}<16'b0100010011010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100010011010100) && ({row_reg, col_reg}<16'b0100010011010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010011010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010011011000) && ({row_reg, col_reg}<16'b0100010011011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010011011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100010011011101) && ({row_reg, col_reg}<16'b0100010011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010011011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100010011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010011100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010011100010) && ({row_reg, col_reg}<16'b0100010011100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010011100100) && ({row_reg, col_reg}<16'b0100010011100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010011100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010011100111) && ({row_reg, col_reg}<16'b0100010011101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010011101010) && ({row_reg, col_reg}<16'b0100010011101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100010011101101) && ({row_reg, col_reg}<16'b0100010011110001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0100010011110001) && ({row_reg, col_reg}<16'b0100010100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010100000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010100000001) && ({row_reg, col_reg}<16'b0100010100000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010100000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100010100000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100010100000101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100010100000110)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100010100000111) && ({row_reg, col_reg}<16'b0100010100001001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100010100001001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100010100001010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100010100001011)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100010100001100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100010100001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100010100001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100010100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010100010000) && ({row_reg, col_reg}<16'b0100010100010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010100010011) && ({row_reg, col_reg}<16'b0100010100010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010100010101) && ({row_reg, col_reg}<16'b0100010100011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100010100011001) && ({row_reg, col_reg}<16'b0100010100011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100010100011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100010100011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010100011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010100011111) && ({row_reg, col_reg}<16'b0100010100100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100010100100001) && ({row_reg, col_reg}<16'b0100010100100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100010100100100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100010100100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100010100100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100010100100111) && ({row_reg, col_reg}<16'b0100010100101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010100101011) && ({row_reg, col_reg}<16'b0100010100101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100010100101101) && ({row_reg, col_reg}<16'b0100010100110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100010100110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100010100110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100010100110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100010100110011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==16'b0100010100110100)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100010100110101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100010100110110)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0100010100110111) && ({row_reg, col_reg}<16'b0100010100111001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100010100111001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100010100111010) && ({row_reg, col_reg}<16'b0100010100111101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100010100111101)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100010100111110) && ({row_reg, col_reg}<16'b0100010101000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100010101000000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100010101000001)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0100010101000010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0100010101000011) && ({row_reg, col_reg}<16'b0100010101000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100010101000110) && ({row_reg, col_reg}<16'b0100010101001001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100010101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100010101001010) && ({row_reg, col_reg}<16'b0100010101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010101001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100010101001101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100010101001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100010101001111) && ({row_reg, col_reg}<16'b0100010101010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100010101010011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0100010101010100) && ({row_reg, col_reg}<16'b0100010101011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010101011001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0100010101011010) && ({row_reg, col_reg}<16'b0100010101011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100010101011111) && ({row_reg, col_reg}<16'b0100010101100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100010101100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100010101100011) && ({row_reg, col_reg}<16'b0100010101100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010101100101) && ({row_reg, col_reg}<16'b0100010101100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100010101100111) && ({row_reg, col_reg}<16'b0100010101101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100010101101001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100010101101010) && ({row_reg, col_reg}<16'b0100010101101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010101101100) && ({row_reg, col_reg}<16'b0100010101101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100010101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010101101111) && ({row_reg, col_reg}<16'b0100010101110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010101110011) && ({row_reg, col_reg}<16'b0100010101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010101110110) && ({row_reg, col_reg}<16'b0100010101111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010101111101) && ({row_reg, col_reg}<16'b0100010101111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010101111111) && ({row_reg, col_reg}<16'b0100010110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010110000011) && ({row_reg, col_reg}<16'b0100010110100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010110100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100010110100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010110100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010110100101) && ({row_reg, col_reg}<16'b0100010110101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010110101100) && ({row_reg, col_reg}<16'b0100010110101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010110101110) && ({row_reg, col_reg}<16'b0100010110110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010110110001) && ({row_reg, col_reg}<16'b0100010110110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010110110100) && ({row_reg, col_reg}<16'b0100010110110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010110110110) && ({row_reg, col_reg}<16'b0100010110111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010110111000) && ({row_reg, col_reg}<16'b0100010110111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010110111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100010110111011) && ({row_reg, col_reg}<16'b0100010110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010110111110) && ({row_reg, col_reg}<16'b0100010111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010111000000) && ({row_reg, col_reg}<16'b0100010111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100010111000011) && ({row_reg, col_reg}<16'b0100010111000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010111000101) && ({row_reg, col_reg}<16'b0100010111001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010111001010) && ({row_reg, col_reg}<16'b0100010111010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100010111010100) && ({row_reg, col_reg}<16'b0100010111011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010111011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100010111011101) && ({row_reg, col_reg}<16'b0100010111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010111011111) && ({row_reg, col_reg}<16'b0100010111100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010111100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010111100010) && ({row_reg, col_reg}<16'b0100010111100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010111100111) && ({row_reg, col_reg}<16'b0100010111101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010111101001) && ({row_reg, col_reg}<16'b0100010111110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100010111110000)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0100010111110001) && ({row_reg, col_reg}<16'b0100011000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100011000000000) && ({row_reg, col_reg}<16'b0100011000000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011000000011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100011000000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100011000000101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100011000000110)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}>=16'b0100011000000111) && ({row_reg, col_reg}<16'b0100011000001001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100011000001001) && ({row_reg, col_reg}<16'b0100011000001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100011000001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011000001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100011000001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011000010000) && ({row_reg, col_reg}<16'b0100011000010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100011000010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011000010011) && ({row_reg, col_reg}<16'b0100011000010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011000010101) && ({row_reg, col_reg}<16'b0100011000011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100011000011001) && ({row_reg, col_reg}<16'b0100011000011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100011000011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100011000011101) && ({row_reg, col_reg}<16'b0100011000100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100011000100010) && ({row_reg, col_reg}<16'b0100011000100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100011000100100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100011000100101) && ({row_reg, col_reg}<16'b0100011000100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011000100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100011000101000) && ({row_reg, col_reg}<16'b0100011000101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011000101011) && ({row_reg, col_reg}<16'b0100011000101110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100011000101110) && ({row_reg, col_reg}<16'b0100011000110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100011000110000) && ({row_reg, col_reg}<16'b0100011000110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100011000110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011000110011)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0100011000110100) && ({row_reg, col_reg}<16'b0100011000110111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100011000110111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0100011000111000) && ({row_reg, col_reg}<16'b0100011000111010)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0100011000111010) && ({row_reg, col_reg}<16'b0100011000111100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100011000111100) && ({row_reg, col_reg}<16'b0100011001000000)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100011001000000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100011001000001)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100011001000010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0100011001000011) && ({row_reg, col_reg}<16'b0100011001000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100011001000110) && ({row_reg, col_reg}<16'b0100011001001001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100011001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100011001001010) && ({row_reg, col_reg}<16'b0100011001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100011001001100) && ({row_reg, col_reg}<16'b0100011001001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100011001001111) && ({row_reg, col_reg}<16'b0100011001010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011001010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100011001010100) && ({row_reg, col_reg}<16'b0100011001010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011001010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011001010111) && ({row_reg, col_reg}<16'b0100011001011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011001011001)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0100011001011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100011001011011) && ({row_reg, col_reg}<16'b0100011001011101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100011001011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100011001011110) && ({row_reg, col_reg}<16'b0100011001100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100011001100000) && ({row_reg, col_reg}<16'b0100011001100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100011001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100011001100011) && ({row_reg, col_reg}<16'b0100011001101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100011001101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100011001101001) && ({row_reg, col_reg}<16'b0100011001101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011001101100) && ({row_reg, col_reg}<16'b0100011001101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100011001101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011001110000) && ({row_reg, col_reg}<16'b0100011001110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011001110010) && ({row_reg, col_reg}<16'b0100011001110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011001110110) && ({row_reg, col_reg}<16'b0100011001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011010000000) && ({row_reg, col_reg}<16'b0100011010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011010000011) && ({row_reg, col_reg}<16'b0100011010100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100011010100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100011010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011010100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100011010100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011010100110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011010100111) && ({row_reg, col_reg}<16'b0100011010101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011010101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011010101101) && ({row_reg, col_reg}<16'b0100011010110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011010110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100011010110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011010110110) && ({row_reg, col_reg}<16'b0100011010111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011010111000) && ({row_reg, col_reg}<16'b0100011010111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011010111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100011010111011) && ({row_reg, col_reg}<16'b0100011010111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011010111101) && ({row_reg, col_reg}<16'b0100011010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100011010111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011011000000) && ({row_reg, col_reg}<16'b0100011011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100011011000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011011000100) && ({row_reg, col_reg}<16'b0100011011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011011001001) && ({row_reg, col_reg}<16'b0100011011001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100011011001011) && ({row_reg, col_reg}<16'b0100011011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011011001110) && ({row_reg, col_reg}<16'b0100011011010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100011011010001) && ({row_reg, col_reg}<16'b0100011011010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011011010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100011011010100) && ({row_reg, col_reg}<16'b0100011011010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011011010111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100011011011000) && ({row_reg, col_reg}<16'b0100011011011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011011011100) && ({row_reg, col_reg}<16'b0100011011011110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100011011011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011011011111) && ({row_reg, col_reg}<16'b0100011011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100011011100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011011100010) && ({row_reg, col_reg}<16'b0100011011100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011011100101) && ({row_reg, col_reg}<16'b0100011011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011011100111) && ({row_reg, col_reg}<16'b0100011011101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011011101001) && ({row_reg, col_reg}<16'b0100011011101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100011011101111) && ({row_reg, col_reg}<16'b0100011011110001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0100011011110001) && ({row_reg, col_reg}<16'b0100011100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100011100000000) && ({row_reg, col_reg}<16'b0100011100000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011100000011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100011100000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100011100000101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0100011100000110) && ({row_reg, col_reg}<16'b0100011100001000)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0100011100001000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100011100001001) && ({row_reg, col_reg}<16'b0100011100001011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100011100001011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011100001100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0100011100001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011100001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100011100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011100010000) && ({row_reg, col_reg}<16'b0100011100010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100011100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011100010011) && ({row_reg, col_reg}<16'b0100011100010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011100010101) && ({row_reg, col_reg}<16'b0100011100011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100011100011001) && ({row_reg, col_reg}<16'b0100011100011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100011100011100) && ({row_reg, col_reg}<16'b0100011100100010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011100100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100011100100011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100011100100100) && ({row_reg, col_reg}<16'b0100011100100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011100100110)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0100011100100111) && ({row_reg, col_reg}<16'b0100011100101001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100011100101001) && ({row_reg, col_reg}<16'b0100011100101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100011100101011) && ({row_reg, col_reg}<16'b0100011100110011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011100110011)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0100011100110100) && ({row_reg, col_reg}<16'b0100011100111000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011100111000)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0100011100111001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100011100111010)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100011100111011) && ({row_reg, col_reg}<16'b0100011100111101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100011100111101)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100011100111110) && ({row_reg, col_reg}<16'b0100011101000010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100011101000010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100011101000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011101000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011101000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100011101000110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0100011101000111) && ({row_reg, col_reg}<16'b0100011101001001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100011101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100011101001010) && ({row_reg, col_reg}<16'b0100011101001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011101001100) && ({row_reg, col_reg}<16'b0100011101001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100011101001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100011101001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100011101010000) && ({row_reg, col_reg}<16'b0100011101010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100011101010011) && ({row_reg, col_reg}<16'b0100011101010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100011101010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100011101010110) && ({row_reg, col_reg}<16'b0100011101011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011101011000) && ({row_reg, col_reg}<16'b0100011101011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100011101011010) && ({row_reg, col_reg}<16'b0100011101011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011101011101) && ({row_reg, col_reg}<16'b0100011101100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100011101100011) && ({row_reg, col_reg}<16'b0100011101100110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100011101100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011101100111) && ({row_reg, col_reg}<16'b0100011101101001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100011101101001) && ({row_reg, col_reg}<16'b0100011101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100011101101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011101101101) && ({row_reg, col_reg}<16'b0100011101110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100011101110000) && ({row_reg, col_reg}<16'b0100011101110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011101110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100011101110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100011101110100) && ({row_reg, col_reg}<16'b0100011101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011101110110) && ({row_reg, col_reg}<16'b0100011101111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011101111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100011101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011101111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011101111101) && ({row_reg, col_reg}<16'b0100011110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011110000000) && ({row_reg, col_reg}<16'b0100011110000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011110000010) && ({row_reg, col_reg}<16'b0100011110100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100011110100001) && ({row_reg, col_reg}<16'b0100011110100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100011110100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011110100100) && ({row_reg, col_reg}<16'b0100011110100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011110100110) && ({row_reg, col_reg}<16'b0100011110101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011110101000) && ({row_reg, col_reg}<16'b0100011110101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011110101011) && ({row_reg, col_reg}<16'b0100011110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011110101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011110101110) && ({row_reg, col_reg}<16'b0100011110110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011110110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011110110010) && ({row_reg, col_reg}<16'b0100011110110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011110110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100011110110101) && ({row_reg, col_reg}<16'b0100011110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011110111101) && ({row_reg, col_reg}<16'b0100011111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011111000000) && ({row_reg, col_reg}<16'b0100011111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100011111000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011111000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011111000101) && ({row_reg, col_reg}<16'b0100011111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011111001001) && ({row_reg, col_reg}<16'b0100011111001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100011111001011) && ({row_reg, col_reg}<16'b0100011111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011111001110) && ({row_reg, col_reg}<16'b0100011111010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100011111010001) && ({row_reg, col_reg}<16'b0100011111011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011111011100) && ({row_reg, col_reg}<16'b0100011111011110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100011111011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011111011111) && ({row_reg, col_reg}<16'b0100011111100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100011111100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011111100010) && ({row_reg, col_reg}<16'b0100011111100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011111100110) && ({row_reg, col_reg}<16'b0100011111101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100011111101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011111101001) && ({row_reg, col_reg}<16'b0100011111101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100011111101101) && ({row_reg, col_reg}<16'b0100011111110001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0100011111110001) && ({row_reg, col_reg}<16'b0100100000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100100000000000) && ({row_reg, col_reg}<16'b0100100000000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100100000000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100100000000011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100100000000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0100100000000101) && ({row_reg, col_reg}<16'b0100100000001011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100100000001011) && ({row_reg, col_reg}<16'b0100100000001101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0100100000001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100000001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100100000001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100000010000) && ({row_reg, col_reg}<16'b0100100000010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100100000010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100000010011) && ({row_reg, col_reg}<16'b0100100000010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100000010101) && ({row_reg, col_reg}<16'b0100100000011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100000011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100100000011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100100000011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100100000011100) && ({row_reg, col_reg}<16'b0100100000100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100100000100101) && ({row_reg, col_reg}<16'b0100100000100111)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0100100000100111) && ({row_reg, col_reg}<16'b0100100000110011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100000110011)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0100100000110100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0100100000110101) && ({row_reg, col_reg}<16'b0100100000111000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100000111000)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0100100000111001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100100000111010)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100100000111011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100100000111100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100100000111101)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}>=16'b0100100000111110) && ({row_reg, col_reg}<16'b0100100001000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100001000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100100001000001)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0100100001000010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100001000011)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0100100001000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100100001000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100100001000110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100100001000111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100100001001000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100100001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100100001001010) && ({row_reg, col_reg}<16'b0100100001001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100100001001100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100100001001101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0100100001001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100100001001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100100001010000) && ({row_reg, col_reg}<16'b0100100001010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100100001010010) && ({row_reg, col_reg}<16'b0100100001010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100100001010101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100100001010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100100001010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100001011000) && ({row_reg, col_reg}<16'b0100100001011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100100001011010) && ({row_reg, col_reg}<16'b0100100001100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100001100000) && ({row_reg, col_reg}<16'b0100100001100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100100001100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100100001100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100001100101) && ({row_reg, col_reg}<16'b0100100001100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100100001100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100001101000) && ({row_reg, col_reg}<16'b0100100001101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100001101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100001101110) && ({row_reg, col_reg}<16'b0100100001110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100100001110000) && ({row_reg, col_reg}<16'b0100100001110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100001110010) && ({row_reg, col_reg}<16'b0100100001110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100100001110110) && ({row_reg, col_reg}<16'b0100100001111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100001111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100001111100) && ({row_reg, col_reg}<16'b0100100001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100100001111110) && ({row_reg, col_reg}<16'b0100100010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100010000000) && ({row_reg, col_reg}<16'b0100100010000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100010000010) && ({row_reg, col_reg}<16'b0100100010100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100100010100001) && ({row_reg, col_reg}<16'b0100100010100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100100010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100010100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100010100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100010100110) && ({row_reg, col_reg}<16'b0100100010101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100100010101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100010101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100010101010) && ({row_reg, col_reg}<16'b0100100010110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100010110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100100010110010) && ({row_reg, col_reg}<16'b0100100010110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100010110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100100010110101) && ({row_reg, col_reg}<16'b0100100010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100010111110) && ({row_reg, col_reg}<16'b0100100011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100011000000) && ({row_reg, col_reg}<16'b0100100011000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100100011000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100100011000011) && ({row_reg, col_reg}<16'b0100100011000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100011000101) && ({row_reg, col_reg}<16'b0100100011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100011001000) && ({row_reg, col_reg}<16'b0100100011001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100100011001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100011001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100011001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100011001110) && ({row_reg, col_reg}<16'b0100100011010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100100011010000) && ({row_reg, col_reg}<16'b0100100011011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100011011000) && ({row_reg, col_reg}<16'b0100100011011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100011011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100011011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100100011011101) && ({row_reg, col_reg}<16'b0100100011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100011011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100100011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100100011100001) && ({row_reg, col_reg}<16'b0100100011100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100100011100011) && ({row_reg, col_reg}<16'b0100100011100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100011100101) && ({row_reg, col_reg}<16'b0100100011101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100011101000) && ({row_reg, col_reg}<16'b0100100011101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100011101010) && ({row_reg, col_reg}<16'b0100100011101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100100011101101) && ({row_reg, col_reg}<16'b0100100011110001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0100100011110001) && ({row_reg, col_reg}<16'b0100100100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100100100000000) && ({row_reg, col_reg}<16'b0100100100000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100100100000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100100100000011) && ({row_reg, col_reg}<16'b0100100100000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100100100000101) && ({row_reg, col_reg}<16'b0100100100001000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100100001000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100100100001001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100100100001010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100100100001011) && ({row_reg, col_reg}<16'b0100100100001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100100100001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100100001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100100100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100100100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100100100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100100010011) && ({row_reg, col_reg}<16'b0100100100010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100100010101) && ({row_reg, col_reg}<16'b0100100100011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100100011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100100100011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100100100011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100100011100) && ({row_reg, col_reg}<16'b0100100100100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100100100101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0100100100100110) && ({row_reg, col_reg}<16'b0100100100101001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100100101001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0100100100101010) && ({row_reg, col_reg}<16'b0100100100110001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100100110001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100100100110010) && ({row_reg, col_reg}<16'b0100100100110100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100100110100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100100100110101)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100100100110110) && ({row_reg, col_reg}<16'b0100100100111010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100100100111010)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100100100111011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100100100111100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100100100111101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100100111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100100111111) && ({row_reg, col_reg}<16'b0100100101000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100100101000101) && ({row_reg, col_reg}<16'b0100100101000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100100101000111) && ({row_reg, col_reg}<16'b0100100101001001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100100101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100100101001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100100101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100100101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100100101001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100100101001110) && ({row_reg, col_reg}<16'b0100100101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100100101010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100100101010001) && ({row_reg, col_reg}<16'b0100100101010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100100101010011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100100101010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100100101010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100101010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100100101010111) && ({row_reg, col_reg}<16'b0100100101011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100100101011100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0100100101011101) && ({row_reg, col_reg}<16'b0100100101011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100101011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100100101100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100100101100001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100101100010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100100101100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100100101100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100100101100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100100101100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100101100111) && ({row_reg, col_reg}<16'b0100100101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100101101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100100101101011) && ({row_reg, col_reg}<16'b0100100101101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100101101101) && ({row_reg, col_reg}<16'b0100100101110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100101110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100101110010) && ({row_reg, col_reg}<16'b0100100101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100100101110110) && ({row_reg, col_reg}<16'b0100100101111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100101111100) && ({row_reg, col_reg}<16'b0100100101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100100101111110) && ({row_reg, col_reg}<16'b0100100110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100110000000) && ({row_reg, col_reg}<16'b0100100110000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100110000010) && ({row_reg, col_reg}<16'b0100100110100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100100110100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100100110100011) && ({row_reg, col_reg}<16'b0100100110100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100110100110) && ({row_reg, col_reg}<16'b0100100110101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100100110101000) && ({row_reg, col_reg}<16'b0100100110101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100110101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100110101101) && ({row_reg, col_reg}<16'b0100100110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100110111110) && ({row_reg, col_reg}<16'b0100100111000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100111000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100100111000010) && ({row_reg, col_reg}<16'b0100100111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100111001000) && ({row_reg, col_reg}<16'b0100100111001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100100111001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100111001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100111001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100111001110) && ({row_reg, col_reg}<16'b0100100111010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100100111010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100111010001) && ({row_reg, col_reg}<16'b0100100111010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100100111010100) && ({row_reg, col_reg}<16'b0100100111010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100111010111) && ({row_reg, col_reg}<16'b0100100111011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100111011010) && ({row_reg, col_reg}<16'b0100100111011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100111011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100100111011101) && ({row_reg, col_reg}<16'b0100100111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100111011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100100111100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100100111100001) && ({row_reg, col_reg}<16'b0100100111100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100100111100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100111100100) && ({row_reg, col_reg}<16'b0100100111100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100111100111) && ({row_reg, col_reg}<16'b0100100111101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100111101010) && ({row_reg, col_reg}<16'b0100100111101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100100111101111) && ({row_reg, col_reg}<16'b0100100111110001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0100100111110001) && ({row_reg, col_reg}<16'b0100101000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100101000000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100101000000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101000000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100101000000011) && ({row_reg, col_reg}<16'b0100101000000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100101000000101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100101000000110)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}>=16'b0100101000000111) && ({row_reg, col_reg}<16'b0100101000001001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100101000001001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100101000001010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100101000001011)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100101000001100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100101000001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100101000001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101000001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100101000010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100101000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100101000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101000010011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100101000010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101000010101) && ({row_reg, col_reg}<16'b0100101000011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100101000011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100101000011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101000011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100101000011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101000011100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100101000011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100101000011110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100101000011111) && ({row_reg, col_reg}<16'b0100101000100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101000100101) && ({row_reg, col_reg}<16'b0100101000101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100101000101010) && ({row_reg, col_reg}<16'b0100101000110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101000110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100101000110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101000110011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100101000110100) && ({row_reg, col_reg}<16'b0100101000111000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100101000111000) && ({row_reg, col_reg}<16'b0100101000111010)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100101000111010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100101000111011)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100101000111100) && ({row_reg, col_reg}<16'b0100101000111110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100101000111110) && ({row_reg, col_reg}<16'b0100101001000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100101001000000) && ({row_reg, col_reg}<16'b0100101001000010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100101001000010) && ({row_reg, col_reg}<16'b0100101001000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100101001000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101001000101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100101001000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100101001000111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100101001001000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100101001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100101001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101001001100) && ({row_reg, col_reg}<16'b0100101001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101001010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100101001010001) && ({row_reg, col_reg}<16'b0100101001010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100101001010100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0100101001010101) && ({row_reg, col_reg}<16'b0100101001010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100101001010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100101001011000) && ({row_reg, col_reg}<16'b0100101001011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100101001011100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0100101001011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100101001011110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0100101001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101001100000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0100101001100001) && ({row_reg, col_reg}<16'b0100101001100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100101001100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101001100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100101001100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101001100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101001100111) && ({row_reg, col_reg}<16'b0100101001101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100101001101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101001101101) && ({row_reg, col_reg}<16'b0100101001110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101001110001) && ({row_reg, col_reg}<16'b0100101001110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101001110011) && ({row_reg, col_reg}<16'b0100101001110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101001110110) && ({row_reg, col_reg}<16'b0100101001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101001111011) && ({row_reg, col_reg}<16'b0100101001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100101001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101010000000) && ({row_reg, col_reg}<16'b0100101010000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101010000010) && ({row_reg, col_reg}<16'b0100101010100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100101010100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101010100011) && ({row_reg, col_reg}<16'b0100101010100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101010100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101010100110) && ({row_reg, col_reg}<16'b0100101010101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101010101000) && ({row_reg, col_reg}<16'b0100101010101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101010101011) && ({row_reg, col_reg}<16'b0100101010101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101010101101) && ({row_reg, col_reg}<16'b0100101010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101010110110) && ({row_reg, col_reg}<16'b0100101010111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101010111000) && ({row_reg, col_reg}<16'b0100101010111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101010111111) && ({row_reg, col_reg}<16'b0100101011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101011000001) && ({row_reg, col_reg}<16'b0100101011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101011001110) && ({row_reg, col_reg}<16'b0100101011010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100101011010100) && ({row_reg, col_reg}<16'b0100101011010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101011010111) && ({row_reg, col_reg}<16'b0100101011011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101011011001) && ({row_reg, col_reg}<16'b0100101011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101011011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100101011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101011100001) && ({row_reg, col_reg}<16'b0100101011100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101011100011) && ({row_reg, col_reg}<16'b0100101011100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101011100101) && ({row_reg, col_reg}<16'b0100101011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101011100111) && ({row_reg, col_reg}<16'b0100101011101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101011101001) && ({row_reg, col_reg}<16'b0100101011110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100101011110000)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0100101011110001) && ({row_reg, col_reg}<16'b0100101100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100101100000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100101100000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101100000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101100000011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100101100000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100101100000101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100101100000110)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}>=16'b0100101100000111) && ({row_reg, col_reg}<16'b0100101100001010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100101100001010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100101100001011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100101100001100)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0100101100001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100101100001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101100010000) && ({row_reg, col_reg}<16'b0100101100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100101100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101100010011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100101100010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101100010101) && ({row_reg, col_reg}<16'b0100101100011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100101100011000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100101100011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100101100011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101100011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100101100011100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100101100011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101100011110) && ({row_reg, col_reg}<16'b0100101100100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100101100100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100101100101000) && ({row_reg, col_reg}<16'b0100101100101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100101100101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101100101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100101100110000) && ({row_reg, col_reg}<16'b0100101100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100101100110011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100101100110100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100101100110101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100101100110110) && ({row_reg, col_reg}<16'b0100101100111010)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100101100111010) && ({row_reg, col_reg}<16'b0100101100111100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100101100111100)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0100101100111101) && ({row_reg, col_reg}<16'b0100101101000010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100101101000010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100101101000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100101101000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101101000101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100101101000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100101101000111) && ({row_reg, col_reg}<16'b0100101101001001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100101101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100101101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101101001100) && ({row_reg, col_reg}<16'b0100101101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100101101010000) && ({row_reg, col_reg}<16'b0100101101010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100101101010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100101101010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100101101010101)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0100101101010110) && ({row_reg, col_reg}<16'b0100101101011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100101101011000) && ({row_reg, col_reg}<16'b0100101101011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100101101011100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0100101101011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100101101011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0100101101011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101101100000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0100101101100001) && ({row_reg, col_reg}<16'b0100101101100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100101101100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100101101100100) && ({row_reg, col_reg}<16'b0100101101100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101101100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101101100111) && ({row_reg, col_reg}<16'b0100101101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100101101101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101101101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101101101110) && ({row_reg, col_reg}<16'b0100101101110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100101101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101101110001) && ({row_reg, col_reg}<16'b0100101101110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100101101110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101101110100) && ({row_reg, col_reg}<16'b0100101101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101101110110) && ({row_reg, col_reg}<16'b0100101101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101101111000) && ({row_reg, col_reg}<16'b0100101101111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100101101111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101101111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100101101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101101111101) && ({row_reg, col_reg}<16'b0100101110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101110000000) && ({row_reg, col_reg}<16'b0100101110000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101110000010) && ({row_reg, col_reg}<16'b0100101110100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100101110100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101110100011) && ({row_reg, col_reg}<16'b0100101110100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101110100110) && ({row_reg, col_reg}<16'b0100101110101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101110101000) && ({row_reg, col_reg}<16'b0100101110110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101110110001) && ({row_reg, col_reg}<16'b0100101110110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101110110111) && ({row_reg, col_reg}<16'b0100101110111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101110111001) && ({row_reg, col_reg}<16'b0100101111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101111000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100101111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101111000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101111000011) && ({row_reg, col_reg}<16'b0100101111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101111000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101111000110) && ({row_reg, col_reg}<16'b0100101111001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101111001100) && ({row_reg, col_reg}<16'b0100101111010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100101111010100) && ({row_reg, col_reg}<16'b0100101111010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101111010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101111011000) && ({row_reg, col_reg}<16'b0100101111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101111011111) && ({row_reg, col_reg}<16'b0100101111100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101111100001) && ({row_reg, col_reg}<16'b0100101111100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101111100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101111100111) && ({row_reg, col_reg}<16'b0100101111101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101111101001) && ({row_reg, col_reg}<16'b0100101111101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100101111101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101111101101) && ({row_reg, col_reg}<16'b0100101111110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100101111110000)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0100101111110001) && ({row_reg, col_reg}<16'b0100110000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100110000000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100110000000001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0100110000000010) && ({row_reg, col_reg}<16'b0100110000000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100110000000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100110000000101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100110000000110)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0100110000000111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100110000001000)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100110000001001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100110000001010)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0100110000001011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100110000001100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100110000001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100110000001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110000001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100110000010000) && ({row_reg, col_reg}<16'b0100110000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100110000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110000010011) && ({row_reg, col_reg}<16'b0100110000010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110000010101)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0100110000010110) && ({row_reg, col_reg}<16'b0100110000011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100110000011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100110000011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110000011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100110000011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100110000011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100110000011110) && ({row_reg, col_reg}<16'b0100110000100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100110000100111) && ({row_reg, col_reg}<16'b0100110000101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100110000101001) && ({row_reg, col_reg}<16'b0100110000101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100110000101110) && ({row_reg, col_reg}<16'b0100110000110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100110000110000) && ({row_reg, col_reg}<16'b0100110000110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110000110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100110000110011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100110000110100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100110000110101)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100110000110110) && ({row_reg, col_reg}<16'b0100110000111001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100110000111001)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0100110000111010)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100110000111011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100110000111100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100110000111101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100110000111110)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0100110000111111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100110001000000)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0100110001000001)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==16'b0100110001000010)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100110001000011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100110001000100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100110001000101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100110001000110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0100110001000111) && ({row_reg, col_reg}<16'b0100110001001001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100110001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100110001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100110001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100110001001100) && ({row_reg, col_reg}<16'b0100110001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100110001010000) && ({row_reg, col_reg}<16'b0100110001010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100110001010011) && ({row_reg, col_reg}<16'b0100110001010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100110001010110) && ({row_reg, col_reg}<16'b0100110001011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100110001011001) && ({row_reg, col_reg}<16'b0100110001011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100110001011100) && ({row_reg, col_reg}<16'b0100110001011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100110001011111) && ({row_reg, col_reg}<16'b0100110001100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100110001100011) && ({row_reg, col_reg}<16'b0100110001100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100110001100110) && ({row_reg, col_reg}<16'b0100110001101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100110001101000) && ({row_reg, col_reg}<16'b0100110001101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110001101100) && ({row_reg, col_reg}<16'b0100110001101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110001101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110001101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100110001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110001110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110001110010) && ({row_reg, col_reg}<16'b0100110001110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110001110100) && ({row_reg, col_reg}<16'b0100110001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110001111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100110001111001) && ({row_reg, col_reg}<16'b0100110001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110001111011) && ({row_reg, col_reg}<16'b0100110001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100110001111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110010000000) && ({row_reg, col_reg}<16'b0100110010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110010000011) && ({row_reg, col_reg}<16'b0100110010100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100110010100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110010100011) && ({row_reg, col_reg}<16'b0100110010100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110010100110) && ({row_reg, col_reg}<16'b0100110010101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100110010101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100110010101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110010101010) && ({row_reg, col_reg}<16'b0100110010110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100110010110001) && ({row_reg, col_reg}<16'b0100110010110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110010110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110010110111) && ({row_reg, col_reg}<16'b0100110010111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110010111001) && ({row_reg, col_reg}<16'b0100110011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110011000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110011000010) && ({row_reg, col_reg}<16'b0100110011000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110011000101) && ({row_reg, col_reg}<16'b0100110011001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110011001000) && ({row_reg, col_reg}<16'b0100110011001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110011001011) && ({row_reg, col_reg}<16'b0100110011010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100110011010011) && ({row_reg, col_reg}<16'b0100110011011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110011011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110011011010) && ({row_reg, col_reg}<16'b0100110011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110011011111) && ({row_reg, col_reg}<16'b0100110011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110011100001) && ({row_reg, col_reg}<16'b0100110011101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110011101001) && ({row_reg, col_reg}<16'b0100110011101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100110011101100) && ({row_reg, col_reg}<16'b0100110011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110011101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100110011110000)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0100110011110001) && ({row_reg, col_reg}<16'b0100110100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100110100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110100000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100110100000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110100000011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0100110100000100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0100110100000101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100110100000110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100110100000111) && ({row_reg, col_reg}<16'b0100110100001010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100110100001010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100110100001011) && ({row_reg, col_reg}<16'b0100110100001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100110100001101) && ({row_reg, col_reg}<16'b0100110100001111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100110100001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100110100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110100010001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100110100010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100110100010011) && ({row_reg, col_reg}<16'b0100110100010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100110100010110) && ({row_reg, col_reg}<16'b0100110100011001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0100110100011001) && ({row_reg, col_reg}<16'b0100110100011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100110100011100) && ({row_reg, col_reg}<16'b0100110100100101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0100110100100101) && ({row_reg, col_reg}<16'b0100110100100111)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0100110100100111) && ({row_reg, col_reg}<16'b0100110100101011)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0100110100101011) && ({row_reg, col_reg}<16'b0100110100101101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0100110100101101) && ({row_reg, col_reg}<16'b0100110100101111)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0100110100101111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100110100110000)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0100110100110001) && ({row_reg, col_reg}<16'b0100110100110011)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0100110100110011) && ({row_reg, col_reg}<16'b0100110100110101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100110100110101) && ({row_reg, col_reg}<16'b0100110100110111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100110100110111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100110100111000) && ({row_reg, col_reg}<16'b0100110100111010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100110100111010)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0100110100111011) && ({row_reg, col_reg}<16'b0100110101000010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100110101000010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100110101000011)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100110101000100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100110101000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100110101000110) && ({row_reg, col_reg}<16'b0100110101001001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100110101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100110101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100110101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100110101001101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0100110101001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100110101001111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0100110101010000) && ({row_reg, col_reg}<16'b0100110101010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100110101010011) && ({row_reg, col_reg}<16'b0100110101010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100110101010110) && ({row_reg, col_reg}<16'b0100110101011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100110101011001) && ({row_reg, col_reg}<16'b0100110101011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100110101011011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0100110101011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100110101011101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100110101011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100110101011111) && ({row_reg, col_reg}<16'b0100110101100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100110101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110101100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100110101100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100110101100101) && ({row_reg, col_reg}<16'b0100110101100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100110101100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100110101101000) && ({row_reg, col_reg}<16'b0100110101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100110101101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110101101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100110101101110) && ({row_reg, col_reg}<16'b0100110101110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100110101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110101110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110101110010) && ({row_reg, col_reg}<16'b0100110101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110101110100) && ({row_reg, col_reg}<16'b0100110101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110101111011) && ({row_reg, col_reg}<16'b0100110101111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110101111101) && ({row_reg, col_reg}<16'b0100110101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110110000000) && ({row_reg, col_reg}<16'b0100110110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110110000011) && ({row_reg, col_reg}<16'b0100110110100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100110110100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100110110100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110110100100) && ({row_reg, col_reg}<16'b0100110110100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110110100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110110100111) && ({row_reg, col_reg}<16'b0100110110101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110110101011) && ({row_reg, col_reg}<16'b0100110110110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100110110110001) && ({row_reg, col_reg}<16'b0100110110110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110110110011) && ({row_reg, col_reg}<16'b0100110110110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110110110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110110110111) && ({row_reg, col_reg}<16'b0100110110111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110110111010) && ({row_reg, col_reg}<16'b0100110111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110111000000) && ({row_reg, col_reg}<16'b0100110111000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110111000011) && ({row_reg, col_reg}<16'b0100110111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110111000111) && ({row_reg, col_reg}<16'b0100110111001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110111001001) && ({row_reg, col_reg}<16'b0100110111001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110111001100) && ({row_reg, col_reg}<16'b0100110111010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100110111010000) && ({row_reg, col_reg}<16'b0100110111011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110111011000) && ({row_reg, col_reg}<16'b0100110111011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110111011010) && ({row_reg, col_reg}<16'b0100110111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110111011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100110111100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110111100001) && ({row_reg, col_reg}<16'b0100110111100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110111100110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110111100111) && ({row_reg, col_reg}<16'b0100110111101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110111101010) && ({row_reg, col_reg}<16'b0100110111101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100110111101101) && ({row_reg, col_reg}<16'b0100110111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110111101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100110111110000)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0100110111110001) && ({row_reg, col_reg}<16'b0100111000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100111000000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100111000000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111000000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111000000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100111000000100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100111000000101) && ({row_reg, col_reg}<16'b0100111000000111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100111000000111) && ({row_reg, col_reg}<16'b0100111000001010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100111000001010) && ({row_reg, col_reg}<16'b0100111000001100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100111000001100) && ({row_reg, col_reg}<16'b0100111000001111)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100111000001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100111000010000)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0100111000010001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100111000010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100111000010011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100111000010100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0100111000010101) && ({row_reg, col_reg}<16'b0100111000011001)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0100111000011001) && ({row_reg, col_reg}<16'b0100111000011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0100111000011011) && ({row_reg, col_reg}<16'b0100111000011101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0100111000011101) && ({row_reg, col_reg}<16'b0100111000011111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100111000011111)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100111000100000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0100111000100001) && ({row_reg, col_reg}<16'b0100111000100101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100111000100101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0100111000100110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100111000100111)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100111000101000)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100111000101001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100111000101010)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0100111000101011) && ({row_reg, col_reg}<16'b0100111000101101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100111000101101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0100111000101110) && ({row_reg, col_reg}<16'b0100111000110000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100111000110000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0100111000110001) && ({row_reg, col_reg}<16'b0100111000110011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0100111000110011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100111000110100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100111000110101)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}>=16'b0100111000110110) && ({row_reg, col_reg}<16'b0100111000111001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100111000111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100111000111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100111000111011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100111000111100)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}>=16'b0100111000111101) && ({row_reg, col_reg}<16'b0100111001000011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0100111001000011) && ({row_reg, col_reg}<16'b0100111001000101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100111001000101) && ({row_reg, col_reg}<16'b0100111001000111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0100111001000111)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0100111001001000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100111001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100111001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100111001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100111001001101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0100111001001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100111001001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100111001010000) && ({row_reg, col_reg}<16'b0100111001010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100111001010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100111001010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100111001010101) && ({row_reg, col_reg}<16'b0100111001011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100111001011000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0100111001011001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0100111001011010) && ({row_reg, col_reg}<16'b0100111001011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100111001011100) && ({row_reg, col_reg}<16'b0100111001011111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0100111001011111) && ({row_reg, col_reg}<16'b0100111001100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100111001100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100111001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100111001100011) && ({row_reg, col_reg}<16'b0100111001100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111001100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100111001100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111001100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111001101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111001101001) && ({row_reg, col_reg}<16'b0100111001101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111001101100) && ({row_reg, col_reg}<16'b0100111001101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111001101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100111001101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100111001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111001110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111001110010) && ({row_reg, col_reg}<16'b0100111001110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111001110100) && ({row_reg, col_reg}<16'b0100111001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111001111011) && ({row_reg, col_reg}<16'b0100111001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100111001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100111001111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111010000000) && ({row_reg, col_reg}<16'b0100111010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111010000011) && ({row_reg, col_reg}<16'b0100111010100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100111010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111010100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100111010100101) && ({row_reg, col_reg}<16'b0100111010100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111010100111) && ({row_reg, col_reg}<16'b0100111010101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100111010101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100111010101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111010101011) && ({row_reg, col_reg}<16'b0100111010101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100111010101101) && ({row_reg, col_reg}<16'b0100111010101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111010101111) && ({row_reg, col_reg}<16'b0100111010110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100111010110001) && ({row_reg, col_reg}<16'b0100111010110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111010110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100111010110100) && ({row_reg, col_reg}<16'b0100111010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111010110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111010110111) && ({row_reg, col_reg}<16'b0100111010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100111010111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111010111010) && ({row_reg, col_reg}<16'b0100111011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111011000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111011000001) && ({row_reg, col_reg}<16'b0100111011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111011000011) && ({row_reg, col_reg}<16'b0100111011001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111011001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111011001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111011001110) && ({row_reg, col_reg}<16'b0100111011010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100111011010000) && ({row_reg, col_reg}<16'b0100111011011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111011011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111011011001) && ({row_reg, col_reg}<16'b0100111011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111011011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100111011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111011100001) && ({row_reg, col_reg}<16'b0100111011101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111011101010) && ({row_reg, col_reg}<16'b0100111011101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100111011101101) && ({row_reg, col_reg}<16'b0100111011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111011101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100111011110000)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0100111011110001) && ({row_reg, col_reg}<16'b0100111100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100111100000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111100000010)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}==16'b0100111100000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100111100000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0100111100000101) && ({row_reg, col_reg}<16'b0100111100000111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0100111100000111) && ({row_reg, col_reg}<16'b0100111100001001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100111100001001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100111100001010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100111100001011) && ({row_reg, col_reg}<16'b0100111100001110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100111100001110)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0100111100001111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0100111100010000) && ({row_reg, col_reg}<16'b0100111100010010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100111100010010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100111100010011)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}>=16'b0100111100010100) && ({row_reg, col_reg}<16'b0100111100011011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100111100011011)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==16'b0100111100011100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0100111100011101) && ({row_reg, col_reg}<16'b0100111100011111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0100111100011111) && ({row_reg, col_reg}<16'b0100111100101000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100111100101000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100111100101001)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100111100101010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100111100101011) && ({row_reg, col_reg}<16'b0100111100101110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0100111100101110) && ({row_reg, col_reg}<16'b0100111100110000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100111100110000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100111100110001)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}>=16'b0100111100110010) && ({row_reg, col_reg}<16'b0100111100110100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100111100110100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100111100110101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100111100110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100111100110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111100111000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100111100111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100111100111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100111100111011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0100111100111100) && ({row_reg, col_reg}<16'b0100111101000110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100111101000110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0100111101000111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100111101001000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100111101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100111101001010) && ({row_reg, col_reg}<16'b0100111101001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100111101001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100111101001110) && ({row_reg, col_reg}<16'b0100111101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100111101010000) && ({row_reg, col_reg}<16'b0100111101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100111101010100) && ({row_reg, col_reg}<16'b0100111101011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100111101011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100111101011010) && ({row_reg, col_reg}<16'b0100111101011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0100111101011100) && ({row_reg, col_reg}<16'b0100111101100000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100111101100000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100111101100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100111101100010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100111101100011) && ({row_reg, col_reg}<16'b0100111101100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111101100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100111101101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111101101001) && ({row_reg, col_reg}<16'b0100111101101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100111101101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111101101101) && ({row_reg, col_reg}<16'b0100111101110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100111101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111101110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111101110010) && ({row_reg, col_reg}<16'b0100111101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111101110100) && ({row_reg, col_reg}<16'b0100111101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111101110110) && ({row_reg, col_reg}<16'b0100111101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111101111000) && ({row_reg, col_reg}<16'b0100111101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111101111100) && ({row_reg, col_reg}<16'b0100111110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111110000000) && ({row_reg, col_reg}<16'b0100111110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111110000011) && ({row_reg, col_reg}<16'b0100111110100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100111110100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111110100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111110100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111110100110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111110100111) && ({row_reg, col_reg}<16'b0100111110101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100111110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111110101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100111110101101) && ({row_reg, col_reg}<16'b0100111110110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100111110110001) && ({row_reg, col_reg}<16'b0100111110110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111110110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100111110110100) && ({row_reg, col_reg}<16'b0100111110110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100111110110110) && ({row_reg, col_reg}<16'b0100111110111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100111110111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111110111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111110111100) && ({row_reg, col_reg}<16'b0100111110111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111110111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100111111000000) && ({row_reg, col_reg}<16'b0100111111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111111000011) && ({row_reg, col_reg}<16'b0100111111001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111111001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111111001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111111001110) && ({row_reg, col_reg}<16'b0100111111010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100111111010011) && ({row_reg, col_reg}<16'b0100111111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111111011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100111111100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100111111100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111111100010) && ({row_reg, col_reg}<16'b0100111111100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111111100100) && ({row_reg, col_reg}<16'b0100111111100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100111111100111) && ({row_reg, col_reg}<16'b0100111111101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111111101010) && ({row_reg, col_reg}<16'b0100111111101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100111111101101) && ({row_reg, col_reg}<16'b0100111111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111111101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100111111110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111111110001)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0100111111110010) && ({row_reg, col_reg}<16'b0101000000000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101000000000001) && ({row_reg, col_reg}<16'b0101000000000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000000000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101000000000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101000000000101) && ({row_reg, col_reg}<16'b0101000000000111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101000000000111) && ({row_reg, col_reg}<16'b0101000000001001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101000000001001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0101000000001010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101000000001011) && ({row_reg, col_reg}<16'b0101000000001101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101000000001101)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==16'b0101000000001110)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0101000000001111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101000000010000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101000000010001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101000000010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101000000010011) && ({row_reg, col_reg}<16'b0101000000010110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101000000010110)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0101000000010111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101000000011000) && ({row_reg, col_reg}<16'b0101000000011010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101000000011010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101000000011011) && ({row_reg, col_reg}<16'b0101000000011101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101000000011101) && ({row_reg, col_reg}<16'b0101000000011111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101000000011111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101000000100000)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}>=16'b0101000000100001) && ({row_reg, col_reg}<16'b0101000000100101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101000000100101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101000000100110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101000000100111)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0101000000101000) && ({row_reg, col_reg}<16'b0101000000101011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101000000101011) && ({row_reg, col_reg}<16'b0101000000101101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0101000000101101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101000000101110) && ({row_reg, col_reg}<16'b0101000000110010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101000000110010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101000000110011) && ({row_reg, col_reg}<16'b0101000000110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101000000110101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101000000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000000110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000000111000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101000000111001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101000000111010) && ({row_reg, col_reg}<16'b0101000000111111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101000000111111) && ({row_reg, col_reg}<16'b0101000001000101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101000001000101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101000001000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101000001000111) && ({row_reg, col_reg}<16'b0101000001001001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101000001001001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0101000001001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000001001011) && ({row_reg, col_reg}<16'b0101000001001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000001001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0101000001001110) && ({row_reg, col_reg}<16'b0101000001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101000001010000) && ({row_reg, col_reg}<16'b0101000001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101000001010100) && ({row_reg, col_reg}<16'b0101000001010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000001010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000001011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000001011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101000001011010)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0101000001011011) && ({row_reg, col_reg}<16'b0101000001011101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101000001011101) && ({row_reg, col_reg}<16'b0101000001011111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101000001011111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101000001100000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101000001100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101000001100010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0101000001100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000001100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000001100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101000001100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101000001100111) && ({row_reg, col_reg}<16'b0101000001101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000001101001) && ({row_reg, col_reg}<16'b0101000001101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000001101011) && ({row_reg, col_reg}<16'b0101000001101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000001101101) && ({row_reg, col_reg}<16'b0101000001110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101000001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000001110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000001110010) && ({row_reg, col_reg}<16'b0101000001110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101000001110100) && ({row_reg, col_reg}<16'b0101000001110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000001110110) && ({row_reg, col_reg}<16'b0101000001111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000001111001) && ({row_reg, col_reg}<16'b0101000001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000001111011) && ({row_reg, col_reg}<16'b0101000010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000010000011) && ({row_reg, col_reg}<16'b0101000010100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101000010100100) && ({row_reg, col_reg}<16'b0101000010100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000010100110) && ({row_reg, col_reg}<16'b0101000010101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101000010101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000010101101) && ({row_reg, col_reg}<16'b0101000010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000010110110) && ({row_reg, col_reg}<16'b0101000010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101000010111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000010111001) && ({row_reg, col_reg}<16'b0101000010111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000010111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000010111100) && ({row_reg, col_reg}<16'b0101000010111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000010111111) && ({row_reg, col_reg}<16'b0101000011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000011000001) && ({row_reg, col_reg}<16'b0101000011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101000011000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000011000100) && ({row_reg, col_reg}<16'b0101000011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000011010001) && ({row_reg, col_reg}<16'b0101000011010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101000011010011) && ({row_reg, col_reg}<16'b0101000011011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000011011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000011011001) && ({row_reg, col_reg}<16'b0101000011011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000011011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101000011011101) && ({row_reg, col_reg}<16'b0101000011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000011011111) && ({row_reg, col_reg}<16'b0101000011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101000011100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000011100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000011100011) && ({row_reg, col_reg}<16'b0101000011101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000011101010) && ({row_reg, col_reg}<16'b0101000011101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101000011101101) && ({row_reg, col_reg}<16'b0101000011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000011101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101000011110000)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0101000011110001) && ({row_reg, col_reg}<16'b0101000100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101000100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000100000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000100000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000100000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101000100000100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101000100000101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101000100000110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101000100000111) && ({row_reg, col_reg}<16'b0101000100001001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101000100001001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101000100001010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101000100001011) && ({row_reg, col_reg}<16'b0101000100010000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101000100010000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101000100010001) && ({row_reg, col_reg}<16'b0101000100010011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101000100010011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0101000100010100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101000100010101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0101000100010110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101000100010111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101000100011000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101000100011001) && ({row_reg, col_reg}<16'b0101000100011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101000100011011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101000100011100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101000100011101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0101000100011110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101000100011111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101000100100000) && ({row_reg, col_reg}<16'b0101000100100100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101000100100100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101000100100101)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0101000100100110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101000100100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101000100101000) && ({row_reg, col_reg}<16'b0101000100101010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101000100101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101000100101011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0101000100101100) && ({row_reg, col_reg}<16'b0101000100101110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101000100101110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101000100101111) && ({row_reg, col_reg}<16'b0101000100110001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101000100110001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101000100110010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101000100110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101000100110100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101000100110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101000100110110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101000100110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101000100111000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101000100111001) && ({row_reg, col_reg}<16'b0101000100111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101000100111011) && ({row_reg, col_reg}<16'b0101000100111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101000100111110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0101000100111111) && ({row_reg, col_reg}<16'b0101000101000100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101000101000100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101000101000101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101000101000110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101000101000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000101001000) && ({row_reg, col_reg}<16'b0101000101001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000101001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000101001011) && ({row_reg, col_reg}<16'b0101000101001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000101001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0101000101001110) && ({row_reg, col_reg}<16'b0101000101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101000101010000) && ({row_reg, col_reg}<16'b0101000101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101000101010100) && ({row_reg, col_reg}<16'b0101000101010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101000101010110) && ({row_reg, col_reg}<16'b0101000101011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000101011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101000101011001) && ({row_reg, col_reg}<16'b0101000101011011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101000101011011) && ({row_reg, col_reg}<16'b0101000101100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101000101100000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101000101100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101000101100010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101000101100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000101100100) && ({row_reg, col_reg}<16'b0101000101100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000101100110) && ({row_reg, col_reg}<16'b0101000101101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101000101101000) && ({row_reg, col_reg}<16'b0101000101101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000101101101) && ({row_reg, col_reg}<16'b0101000101110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101000101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000101110001) && ({row_reg, col_reg}<16'b0101000101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101000101110100) && ({row_reg, col_reg}<16'b0101000101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000101110110) && ({row_reg, col_reg}<16'b0101000101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000101111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101000101111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101000101111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000101111011) && ({row_reg, col_reg}<16'b0101000110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000110000011) && ({row_reg, col_reg}<16'b0101000110101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101000110101011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==16'b0101000110101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000110101101) && ({row_reg, col_reg}<16'b0101000110110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000110110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101000110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101000110110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000110111000) && ({row_reg, col_reg}<16'b0101000110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000110111110) && ({row_reg, col_reg}<16'b0101000111000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000111000001) && ({row_reg, col_reg}<16'b0101000111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101000111000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000111000100) && ({row_reg, col_reg}<16'b0101000111000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000111000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101000111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000111001000) && ({row_reg, col_reg}<16'b0101000111001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000111001010) && ({row_reg, col_reg}<16'b0101000111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000111010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101000111010010) && ({row_reg, col_reg}<16'b0101000111010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000111010111) && ({row_reg, col_reg}<16'b0101000111011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000111011010) && ({row_reg, col_reg}<16'b0101000111011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000111011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101000111011101) && ({row_reg, col_reg}<16'b0101000111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000111011111) && ({row_reg, col_reg}<16'b0101000111100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101000111100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000111100010) && ({row_reg, col_reg}<16'b0101000111100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000111100100) && ({row_reg, col_reg}<16'b0101000111101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000111101010) && ({row_reg, col_reg}<16'b0101000111101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101000111101100) && ({row_reg, col_reg}<16'b0101000111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000111101111) && ({row_reg, col_reg}<16'b0101000111110001)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0101000111110001) && ({row_reg, col_reg}<16'b0101001000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101001000000000) && ({row_reg, col_reg}<16'b0101001000000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001000000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101001000000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001000000100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101001000000101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101001000000110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101001000000111) && ({row_reg, col_reg}<16'b0101001000001001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101001000001001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101001000001010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101001000001011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101001000001100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101001000001101) && ({row_reg, col_reg}<16'b0101001000010000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101001000010000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101001000010001) && ({row_reg, col_reg}<16'b0101001000010011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101001000010011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0101001000010100) && ({row_reg, col_reg}<16'b0101001000010110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101001000010110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101001000010111) && ({row_reg, col_reg}<16'b0101001000011001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101001000011001) && ({row_reg, col_reg}<16'b0101001000011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101001000011011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101001000011100) && ({row_reg, col_reg}<16'b0101001000011110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101001000011110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101001000011111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101001000100000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0101001000100001) && ({row_reg, col_reg}<16'b0101001000100011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101001000100011) && ({row_reg, col_reg}<16'b0101001000100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101001000100101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101001000100110) && ({row_reg, col_reg}<16'b0101001000101010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101001000101010) && ({row_reg, col_reg}<16'b0101001000101100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101001000101100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0101001000101101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101001000101110)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101001000101111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101001000110000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101001000110001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101001000110010) && ({row_reg, col_reg}<16'b0101001000110100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101001000110100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101001000110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101001000110110) && ({row_reg, col_reg}<16'b0101001000111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101001000111001) && ({row_reg, col_reg}<16'b0101001000111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101001000111011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0101001000111100) && ({row_reg, col_reg}<16'b0101001000111110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101001000111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101001000111111) && ({row_reg, col_reg}<16'b0101001001000100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101001001000100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101001001000101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101001001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101001001000111) && ({row_reg, col_reg}<16'b0101001001001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001001001001) && ({row_reg, col_reg}<16'b0101001001001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101001001001100) && ({row_reg, col_reg}<16'b0101001001001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101001001001111) && ({row_reg, col_reg}<16'b0101001001010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001001010001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0101001001010010) && ({row_reg, col_reg}<16'b0101001001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101001001010101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0101001001010110) && ({row_reg, col_reg}<16'b0101001001011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101001001011000) && ({row_reg, col_reg}<16'b0101001001011011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001001011011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0101001001011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101001001011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001001011110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0101001001011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001001100000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101001001100001)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0101001001100010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001001100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101001001100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101001001100101) && ({row_reg, col_reg}<16'b0101001001100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101001001100111) && ({row_reg, col_reg}<16'b0101001001101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101001001101001) && ({row_reg, col_reg}<16'b0101001001110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001001110001) && ({row_reg, col_reg}<16'b0101001001110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101001001110100) && ({row_reg, col_reg}<16'b0101001001110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001001110110) && ({row_reg, col_reg}<16'b0101001001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001001111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101001001111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101001001111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101001001111011) && ({row_reg, col_reg}<16'b0101001001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001010000000) && ({row_reg, col_reg}<16'b0101001010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001010000011) && ({row_reg, col_reg}<16'b0101001010100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101001010100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001010100010) && ({row_reg, col_reg}<16'b0101001010101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101001010101011) && ({row_reg, col_reg}<16'b0101001010101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101001010101101) && ({row_reg, col_reg}<16'b0101001010110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001010110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001010110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001010110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001010110110) && ({row_reg, col_reg}<16'b0101001010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101001010111000) && ({row_reg, col_reg}<16'b0101001010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001010111110) && ({row_reg, col_reg}<16'b0101001011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101001011000000) && ({row_reg, col_reg}<16'b0101001011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101001011000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001011000100) && ({row_reg, col_reg}<16'b0101001011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001011001000) && ({row_reg, col_reg}<16'b0101001011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101001011001010) && ({row_reg, col_reg}<16'b0101001011010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001011010101) && ({row_reg, col_reg}<16'b0101001011011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101001011011010) && ({row_reg, col_reg}<16'b0101001011011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001011011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101001011011101) && ({row_reg, col_reg}<16'b0101001011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001011011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101001011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101001011100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001011100010) && ({row_reg, col_reg}<16'b0101001011100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101001011100100) && ({row_reg, col_reg}<16'b0101001011101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001011101010) && ({row_reg, col_reg}<16'b0101001011101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101001011101100) && ({row_reg, col_reg}<16'b0101001011101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001011101110) && ({row_reg, col_reg}<16'b0101001011110001)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0101001011110001) && ({row_reg, col_reg}<16'b0101001100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101001100000000) && ({row_reg, col_reg}<16'b0101001100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001100000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101001100000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101001100000100) && ({row_reg, col_reg}<16'b0101001100000110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101001100000110)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0101001100000111)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101001100001000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101001100001001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0101001100001010) && ({row_reg, col_reg}<16'b0101001100001100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101001100001100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101001100001101) && ({row_reg, col_reg}<16'b0101001100010000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101001100010000) && ({row_reg, col_reg}<16'b0101001100010011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101001100010011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101001100010100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101001100010101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0101001100010110) && ({row_reg, col_reg}<16'b0101001100011001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101001100011001) && ({row_reg, col_reg}<16'b0101001100011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101001100011011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101001100011100) && ({row_reg, col_reg}<16'b0101001100011111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101001100011111) && ({row_reg, col_reg}<16'b0101001100100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101001100100001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101001100100010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101001100100011) && ({row_reg, col_reg}<16'b0101001100100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101001100100101) && ({row_reg, col_reg}<16'b0101001100101010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101001100101010) && ({row_reg, col_reg}<16'b0101001100101100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101001100101100) && ({row_reg, col_reg}<16'b0101001100101110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101001100101110) && ({row_reg, col_reg}<16'b0101001100110000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101001100110000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101001100110001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101001100110010)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0101001100110011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101001100110100) && ({row_reg, col_reg}<16'b0101001100110110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101001100110110)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0101001100110111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0101001100111000) && ({row_reg, col_reg}<16'b0101001100111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101001100111010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001100111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001100111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101001100111101)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}==16'b0101001100111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101001100111111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101001101000000)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}>=16'b0101001101000001) && ({row_reg, col_reg}<16'b0101001101000100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101001101000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101001101000101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101001101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101001101000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001101001000) && ({row_reg, col_reg}<16'b0101001101001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101001101001010) && ({row_reg, col_reg}<16'b0101001101001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001101001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101001101001101) && ({row_reg, col_reg}<16'b0101001101001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101001101001111) && ({row_reg, col_reg}<16'b0101001101010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001101010001)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}>=16'b0101001101010010) && ({row_reg, col_reg}<16'b0101001101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101001101010101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0101001101010110) && ({row_reg, col_reg}<16'b0101001101011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101001101011000) && ({row_reg, col_reg}<16'b0101001101011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101001101011010) && ({row_reg, col_reg}<16'b0101001101011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001101011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001101011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001101011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101001101011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001101100000)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0101001101100001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001101100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101001101100011) && ({row_reg, col_reg}<16'b0101001101100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101001101100101) && ({row_reg, col_reg}<16'b0101001101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101001101101010) && ({row_reg, col_reg}<16'b0101001101101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101001101101101) && ({row_reg, col_reg}<16'b0101001101101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101001101101111) && ({row_reg, col_reg}<16'b0101001101110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001101110001) && ({row_reg, col_reg}<16'b0101001101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101001101110100) && ({row_reg, col_reg}<16'b0101001101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001101110110) && ({row_reg, col_reg}<16'b0101001101111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001101111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101001101111010) && ({row_reg, col_reg}<16'b0101001101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001110000000) && ({row_reg, col_reg}<16'b0101001110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001110000011) && ({row_reg, col_reg}<16'b0101001110100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101001110100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001110100010) && ({row_reg, col_reg}<16'b0101001110101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101001110101011) && ({row_reg, col_reg}<16'b0101001110101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101001110101110) && ({row_reg, col_reg}<16'b0101001110110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001110110011) && ({row_reg, col_reg}<16'b0101001110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001110110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001110110110) && ({row_reg, col_reg}<16'b0101001110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101001110111000) && ({row_reg, col_reg}<16'b0101001110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001110111110) && ({row_reg, col_reg}<16'b0101001111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101001111000000) && ({row_reg, col_reg}<16'b0101001111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101001111000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001111000100) && ({row_reg, col_reg}<16'b0101001111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001111001110) && ({row_reg, col_reg}<16'b0101001111010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101001111010001) && ({row_reg, col_reg}<16'b0101001111010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001111010011) && ({row_reg, col_reg}<16'b0101001111011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101001111011001) && ({row_reg, col_reg}<16'b0101001111011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001111011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101001111011101) && ({row_reg, col_reg}<16'b0101001111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001111011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101001111100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101001111100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101001111100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001111100011) && ({row_reg, col_reg}<16'b0101001111100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101001111100110) && ({row_reg, col_reg}<16'b0101001111101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001111101010) && ({row_reg, col_reg}<16'b0101001111101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101001111101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001111101101) && ({row_reg, col_reg}<16'b0101001111110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001111110000)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0101001111110001) && ({row_reg, col_reg}<16'b0101010000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101010000000000) && ({row_reg, col_reg}<16'b0101010000000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010000000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010000000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101010000000100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101010000000101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101010000000110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101010000000111) && ({row_reg, col_reg}<16'b0101010000001010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101010000001010) && ({row_reg, col_reg}<16'b0101010000001101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101010000001101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010000001110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101010000001111) && ({row_reg, col_reg}<16'b0101010000011001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010000011001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101010000011010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101010000011011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101010000011100) && ({row_reg, col_reg}<16'b0101010000100011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010000100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101010000100100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101010000100101) && ({row_reg, col_reg}<16'b0101010000100111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010000100111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101010000101000) && ({row_reg, col_reg}<16'b0101010000110111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010000110111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101010000111000) && ({row_reg, col_reg}<16'b0101010000111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101010000111010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101010000111011) && ({row_reg, col_reg}<16'b0101010000111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010000111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101010000111111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101010001000000)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}>=16'b0101010001000001) && ({row_reg, col_reg}<16'b0101010001000011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010001000011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101010001000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101010001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101010001000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101010001000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010001001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101010001001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101010001001010) && ({row_reg, col_reg}<16'b0101010001001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010001001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101010001001101) && ({row_reg, col_reg}<16'b0101010001001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101010001001111) && ({row_reg, col_reg}<16'b0101010001010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101010001010001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0101010001010010) && ({row_reg, col_reg}<16'b0101010001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101010001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101010001010101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0101010001010110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101010001010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101010001011000) && ({row_reg, col_reg}<16'b0101010001011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101010001011011) && ({row_reg, col_reg}<16'b0101010001011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010001011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101010001011110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101010001011111) && ({row_reg, col_reg}<16'b0101010001100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101010001100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101010001100011) && ({row_reg, col_reg}<16'b0101010001100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101010001100101) && ({row_reg, col_reg}<16'b0101010001101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010001101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010001101100) && ({row_reg, col_reg}<16'b0101010001101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101010001101110) && ({row_reg, col_reg}<16'b0101010001110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101010001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010001110001) && ({row_reg, col_reg}<16'b0101010001110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101010001110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010001110101) && ({row_reg, col_reg}<16'b0101010010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010010000011) && ({row_reg, col_reg}<16'b0101010010101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101010010101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010010101100) && ({row_reg, col_reg}<16'b0101010010101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010010101110) && ({row_reg, col_reg}<16'b0101010010110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010010110000) && ({row_reg, col_reg}<16'b0101010010110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010010110011) && ({row_reg, col_reg}<16'b0101010010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010010110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010010110110) && ({row_reg, col_reg}<16'b0101010010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101010010111000) && ({row_reg, col_reg}<16'b0101010010111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010010111101) && ({row_reg, col_reg}<16'b0101010011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010011000001) && ({row_reg, col_reg}<16'b0101010011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101010011000011) && ({row_reg, col_reg}<16'b0101010011000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010011000101) && ({row_reg, col_reg}<16'b0101010011001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010011001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010011001101) && ({row_reg, col_reg}<16'b0101010011001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010011001111) && ({row_reg, col_reg}<16'b0101010011010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101010011010001) && ({row_reg, col_reg}<16'b0101010011010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010011010100) && ({row_reg, col_reg}<16'b0101010011010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010011010111) && ({row_reg, col_reg}<16'b0101010011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010011011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101010011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101010011100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010011100010) && ({row_reg, col_reg}<16'b0101010011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010011100111) && ({row_reg, col_reg}<16'b0101010011101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010011101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101010011101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010011101101) && ({row_reg, col_reg}<16'b0101010011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010011110000)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0101010011110001) && ({row_reg, col_reg}<16'b0101010100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101010100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010100000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101010100000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010100000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101010100000100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==16'b0101010100000101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101010100000110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010100000111)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==16'b0101010100001000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010100001001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101010100001010) && ({row_reg, col_reg}<16'b0101010100001100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101010100001100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101010100001101) && ({row_reg, col_reg}<16'b0101010100011001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101010100011001) && ({row_reg, col_reg}<16'b0101010100011011)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0101010100011011)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}>=16'b0101010100011100) && ({row_reg, col_reg}<16'b0101010100100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010100100010)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0101010100100011)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0101010100100100)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0101010100100101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010100100110)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0101010100100111)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0101010100101000)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}>=16'b0101010100101001) && ({row_reg, col_reg}<16'b0101010100110111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010100110111)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0101010100111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101010100111001) && ({row_reg, col_reg}<16'b0101010100111011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101010100111011)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0101010100111100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101010100111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101010100111110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101010100111111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010101000000)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}>=16'b0101010101000001) && ({row_reg, col_reg}<16'b0101010101000011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010101000011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0101010101000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101010101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101010101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010101000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010101001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010101001001) && ({row_reg, col_reg}<16'b0101010101001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101010101001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010101001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101010101001101) && ({row_reg, col_reg}<16'b0101010101001111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0101010101001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101010101010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101010101010001)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0101010101010010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101010101010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101010101010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101010101010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101010101010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010101010111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0101010101011000) && ({row_reg, col_reg}<16'b0101010101011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101010101011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010101011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101010101011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101010101011110) && ({row_reg, col_reg}<16'b0101010101100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101010101100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101010101100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101010101100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101010101100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010101100101) && ({row_reg, col_reg}<16'b0101010101100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101010101100111) && ({row_reg, col_reg}<16'b0101010101101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101010101101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010101101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101010101101101) && ({row_reg, col_reg}<16'b0101010101101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101010101101111) && ({row_reg, col_reg}<16'b0101010101110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010101110001) && ({row_reg, col_reg}<16'b0101010101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101010101110100) && ({row_reg, col_reg}<16'b0101010101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010101110110) && ({row_reg, col_reg}<16'b0101010110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010110000011) && ({row_reg, col_reg}<16'b0101010110101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101010110101100) && ({row_reg, col_reg}<16'b0101010110101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010110101110) && ({row_reg, col_reg}<16'b0101010110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101010110110000) && ({row_reg, col_reg}<16'b0101010110110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010110110010) && ({row_reg, col_reg}<16'b0101010110110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010110110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010110110110) && ({row_reg, col_reg}<16'b0101010110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101010110111000) && ({row_reg, col_reg}<16'b0101010110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010110111101) && ({row_reg, col_reg}<16'b0101010111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010111000001) && ({row_reg, col_reg}<16'b0101010111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101010111000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010111000100) && ({row_reg, col_reg}<16'b0101010111001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010111001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010111001101) && ({row_reg, col_reg}<16'b0101010111001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010111001111) && ({row_reg, col_reg}<16'b0101010111010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101010111010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010111010011) && ({row_reg, col_reg}<16'b0101010111010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010111010110) && ({row_reg, col_reg}<16'b0101010111011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010111011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010111011001) && ({row_reg, col_reg}<16'b0101010111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010111011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101010111100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101010111100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010111100010) && ({row_reg, col_reg}<16'b0101010111100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010111100111) && ({row_reg, col_reg}<16'b0101010111101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010111101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101010111101100) && ({row_reg, col_reg}<16'b0101010111101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010111101110) && ({row_reg, col_reg}<16'b0101010111110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010111110000)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0101010111110001) && ({row_reg, col_reg}<16'b0101011000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011000000000) && ({row_reg, col_reg}<16'b0101011000000010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101011000000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011000000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101011000000100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101011000000101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011000000110)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0101011000000111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011000001000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101011000001001)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0101011000001010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101011000001011)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0101011000001100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101011000001101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101011000001110) && ({row_reg, col_reg}<16'b0101011000010111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011000010111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101011000011000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011000011001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0101011000011010)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0101011000011011)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=16'b0101011000011100) && ({row_reg, col_reg}<16'b0101011000011110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101011000011110) && ({row_reg, col_reg}<16'b0101011000100001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011000100001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101011000100010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0101011000100011)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0101011000100100)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0101011000100101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011000100110)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0101011000100111)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0101011000101000)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0101011000101001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011000101010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101011000101011) && ({row_reg, col_reg}<16'b0101011000111001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011000111001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101011000111010) && ({row_reg, col_reg}<16'b0101011000111100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011000111100)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0101011000111101) && ({row_reg, col_reg}<16'b0101011000111111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101011000111111) && ({row_reg, col_reg}<16'b0101011001000001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011001000001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0101011001000010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101011001000011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011001000100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101011001000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101011001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101011001000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011001001000) && ({row_reg, col_reg}<16'b0101011001001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011001001011) && ({row_reg, col_reg}<16'b0101011001001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011001001101) && ({row_reg, col_reg}<16'b0101011001001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101011001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011001010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101011001010001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101011001010010)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0101011001010011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101011001010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101011001010101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101011001010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101011001010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011001011000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0101011001011001) && ({row_reg, col_reg}<16'b0101011001011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101011001011011) && ({row_reg, col_reg}<16'b0101011001011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101011001011101) && ({row_reg, col_reg}<16'b0101011001100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101011001100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101011001100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101011001100011) && ({row_reg, col_reg}<16'b0101011001100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011001100101) && ({row_reg, col_reg}<16'b0101011001101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101011001101001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101011001101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101011001101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101011001101100) && ({row_reg, col_reg}<16'b0101011001101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101011001101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101011001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011001110001) && ({row_reg, col_reg}<16'b0101011001110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011001110100) && ({row_reg, col_reg}<16'b0101011001110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011001110110) && ({row_reg, col_reg}<16'b0101011001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011001111011) && ({row_reg, col_reg}<16'b0101011010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011010000000) && ({row_reg, col_reg}<16'b0101011010000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101011010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011010000011) && ({row_reg, col_reg}<16'b0101011010101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011010101100) && ({row_reg, col_reg}<16'b0101011010101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101011010101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101011010101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101011010110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011010110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011010110010) && ({row_reg, col_reg}<16'b0101011010110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011010110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011010110110) && ({row_reg, col_reg}<16'b0101011010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011010111000) && ({row_reg, col_reg}<16'b0101011010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011010111110) && ({row_reg, col_reg}<16'b0101011011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011011000000) && ({row_reg, col_reg}<16'b0101011011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101011011000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011011000100) && ({row_reg, col_reg}<16'b0101011011000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011011000110) && ({row_reg, col_reg}<16'b0101011011010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011011010000) && ({row_reg, col_reg}<16'b0101011011010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101011011010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011011010011) && ({row_reg, col_reg}<16'b0101011011010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011011010101) && ({row_reg, col_reg}<16'b0101011011011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011011011000) && ({row_reg, col_reg}<16'b0101011011011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011011011010) && ({row_reg, col_reg}<16'b0101011011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011011011111) && ({row_reg, col_reg}<16'b0101011011100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011011100010) && ({row_reg, col_reg}<16'b0101011011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011011100111) && ({row_reg, col_reg}<16'b0101011011101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011011101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101011011101100) && ({row_reg, col_reg}<16'b0101011011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011011101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101011011110000)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0101011011110001) && ({row_reg, col_reg}<16'b0101011100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011100000000) && ({row_reg, col_reg}<16'b0101011100000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011100000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101011100000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101011100000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101011100000101) && ({row_reg, col_reg}<16'b0101011100000111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011100000111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101011100001000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101011100001001)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0101011100001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011100001011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101011100001100)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0101011100001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101011100001110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101011100001111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011100010000)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}>=16'b0101011100010001) && ({row_reg, col_reg}<16'b0101011100010101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011100010101)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0101011100010110)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}>=16'b0101011100010111) && ({row_reg, col_reg}<16'b0101011100011001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011100011001)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0101011100011010)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==16'b0101011100011011)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=16'b0101011100011100) && ({row_reg, col_reg}<16'b0101011100100000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101011100100000) && ({row_reg, col_reg}<16'b0101011100100010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101011100100010)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0101011100100011)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0101011100100100)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0101011100100101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011100100110)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0101011100100111)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0101011100101000)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}>=16'b0101011100101001) && ({row_reg, col_reg}<16'b0101011100101011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011100101011)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}>=16'b0101011100101100) && ({row_reg, col_reg}<16'b0101011100101110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011100101110)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}>=16'b0101011100101111) && ({row_reg, col_reg}<16'b0101011100111000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101011100111000) && ({row_reg, col_reg}<16'b0101011100111100)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0101011100111100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101011100111101) && ({row_reg, col_reg}<16'b0101011100111111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101011100111111)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0101011101000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101011101000001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101011101000010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101011101000011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101011101000100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0101011101000101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101011101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101011101000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011101001000) && ({row_reg, col_reg}<16'b0101011101001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101011101001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101011101001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011101001101) && ({row_reg, col_reg}<16'b0101011101001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101011101001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101011101010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101011101010001) && ({row_reg, col_reg}<16'b0101011101010100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101011101010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101011101010101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101011101010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101011101010111) && ({row_reg, col_reg}<16'b0101011101011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011101011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101011101011011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0101011101011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101011101011101) && ({row_reg, col_reg}<16'b0101011101011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101011101011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101011101100000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101011101100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101011101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101011101100011) && ({row_reg, col_reg}<16'b0101011101100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011101100101) && ({row_reg, col_reg}<16'b0101011101101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101011101101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101011101101100) && ({row_reg, col_reg}<16'b0101011101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011101101110) && ({row_reg, col_reg}<16'b0101011101110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011101110000) && ({row_reg, col_reg}<16'b0101011101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011101110110) && ({row_reg, col_reg}<16'b0101011101111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101011101111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101011101111001) && ({row_reg, col_reg}<16'b0101011101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011101111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011101111100) && ({row_reg, col_reg}<16'b0101011101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101011101111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011110000000) && ({row_reg, col_reg}<16'b0101011110000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101011110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011110000011) && ({row_reg, col_reg}<16'b0101011110101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011110101100) && ({row_reg, col_reg}<16'b0101011110101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011110101110) && ({row_reg, col_reg}<16'b0101011110110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011110110010) && ({row_reg, col_reg}<16'b0101011110110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011110110110) && ({row_reg, col_reg}<16'b0101011110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011110111000) && ({row_reg, col_reg}<16'b0101011110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011110111110) && ({row_reg, col_reg}<16'b0101011111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011111000000) && ({row_reg, col_reg}<16'b0101011111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011111000011) && ({row_reg, col_reg}<16'b0101011111000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011111000101) && ({row_reg, col_reg}<16'b0101011111001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011111001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011111001100) && ({row_reg, col_reg}<16'b0101011111010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011111010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011111010100) && ({row_reg, col_reg}<16'b0101011111011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011111011000) && ({row_reg, col_reg}<16'b0101011111011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011111011010) && ({row_reg, col_reg}<16'b0101011111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011111011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101011111100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101011111100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011111100010) && ({row_reg, col_reg}<16'b0101011111100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011111100111) && ({row_reg, col_reg}<16'b0101011111101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011111101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101011111101100) && ({row_reg, col_reg}<16'b0101011111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011111101111) && ({row_reg, col_reg}<16'b0101011111110001)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0101011111110001) && ({row_reg, col_reg}<16'b0101100000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101100000000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101100000000001) && ({row_reg, col_reg}<16'b0101100000000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101100000000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101100000000100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101100000000101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0101100000000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101100000000111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101100000001000) && ({row_reg, col_reg}<16'b0101100000001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100000001100)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0101100000001101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0101100000001110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101100000001111)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0101100000010000) && ({row_reg, col_reg}<16'b0101100000010010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101100000010010) && ({row_reg, col_reg}<16'b0101100000010100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101100000010100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101100000010101)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==16'b0101100000010110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101100000010111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101100000011000)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0101100000011001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101100000011010)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0101100000011011) && ({row_reg, col_reg}<16'b0101100000011111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101100000011111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101100000100000) && ({row_reg, col_reg}<16'b0101100000100010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101100000100010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101100000100011)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0101100000100100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101100000100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101100000100110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101100000100111) && ({row_reg, col_reg}<16'b0101100000101001)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}>=16'b0101100000101001) && ({row_reg, col_reg}<16'b0101100000110000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101100000110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101100000110001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0101100000110010) && ({row_reg, col_reg}<16'b0101100000110100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101100000110100) && ({row_reg, col_reg}<16'b0101100000110111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101100000110111) && ({row_reg, col_reg}<16'b0101100000111001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101100000111001)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}>=16'b0101100000111010) && ({row_reg, col_reg}<16'b0101100000111100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101100000111100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101100000111101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101100000111110) && ({row_reg, col_reg}<16'b0101100001000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101100001000011) && ({row_reg, col_reg}<16'b0101100001000101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101100001000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101100001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101100001000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100001001000) && ({row_reg, col_reg}<16'b0101100001001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101100001001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100001001100) && ({row_reg, col_reg}<16'b0101100001001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101100001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100001001111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101100001010000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101100001010001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101100001010010)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0101100001010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101100001010100) && ({row_reg, col_reg}<16'b0101100001010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101100001010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100001011000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101100001011001) && ({row_reg, col_reg}<16'b0101100001011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101100001011011) && ({row_reg, col_reg}<16'b0101100001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101100001100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101100001100011) && ({row_reg, col_reg}<16'b0101100001100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100001100110)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}>=16'b0101100001100111) && ({row_reg, col_reg}<16'b0101100001101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101100001101010) && ({row_reg, col_reg}<16'b0101100001101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100001101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100001101101) && ({row_reg, col_reg}<16'b0101100001110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100001110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100001110001) && ({row_reg, col_reg}<16'b0101100001110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100001110110) && ({row_reg, col_reg}<16'b0101100001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100001111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101100001111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100001111101) && ({row_reg, col_reg}<16'b0101100001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100001111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100010000000) && ({row_reg, col_reg}<16'b0101100010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100010000011) && ({row_reg, col_reg}<16'b0101100010101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100010101001) && ({row_reg, col_reg}<16'b0101100010101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100010101011) && ({row_reg, col_reg}<16'b0101100010110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100010110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100010110010) && ({row_reg, col_reg}<16'b0101100010111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100010111000) && ({row_reg, col_reg}<16'b0101100010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100010111110) && ({row_reg, col_reg}<16'b0101100011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100011000000) && ({row_reg, col_reg}<16'b0101100011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100011000011) && ({row_reg, col_reg}<16'b0101100011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100011001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101100011001111) && ({row_reg, col_reg}<16'b0101100011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100011010001) && ({row_reg, col_reg}<16'b0101100011010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100011010011) && ({row_reg, col_reg}<16'b0101100011010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100011010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100011010110) && ({row_reg, col_reg}<16'b0101100011011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100011011000) && ({row_reg, col_reg}<16'b0101100011011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100011011010) && ({row_reg, col_reg}<16'b0101100011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100011011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101100011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101100011100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100011100010) && ({row_reg, col_reg}<16'b0101100011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100011100111) && ({row_reg, col_reg}<16'b0101100011110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100011110000)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0101100011110001) && ({row_reg, col_reg}<16'b0101100100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100100000000) && ({row_reg, col_reg}<16'b0101100100000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101100100000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101100100000100) && ({row_reg, col_reg}<16'b0101100100000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101100100000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101100100000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100100001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101100100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100100001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101100100001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100100001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101100100001110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101100100001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101100100010000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101100100010001)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0101100100010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101100100010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101100100010100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0101100100010101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0101100100010110) && ({row_reg, col_reg}<16'b0101100100011000)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0101100100011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101100100011001)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0101100100011010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101100100011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101100100011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101100100011101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0101100100011110) && ({row_reg, col_reg}<16'b0101100100100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101100100100000) && ({row_reg, col_reg}<16'b0101100100100010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101100100100010) && ({row_reg, col_reg}<16'b0101100100101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101100100101000)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0101100100101001) && ({row_reg, col_reg}<16'b0101100100101110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101100100101110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101100100101111) && ({row_reg, col_reg}<16'b0101100100110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101100100110010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101100100110011)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0101100100110100) && ({row_reg, col_reg}<16'b0101100100111000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101100100111000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101100100111001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101100100111010)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0101100100111011) && ({row_reg, col_reg}<16'b0101100100111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101100100111110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101100100111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101100101000000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101100101000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101100101000010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0101100101000011) && ({row_reg, col_reg}<16'b0101100101000101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101100101000101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101100101000110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101100101000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100101001000) && ({row_reg, col_reg}<16'b0101100101001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101100101001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101100101001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100101001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101100101001101) && ({row_reg, col_reg}<16'b0101100101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100101001111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101100101010000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101100101010001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0101100101010010) && ({row_reg, col_reg}<16'b0101100101010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101100101010100) && ({row_reg, col_reg}<16'b0101100101010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101100101010110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101100101010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100101011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100101011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100101011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100101011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101100101011100) && ({row_reg, col_reg}<16'b0101100101011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101100101011111) && ({row_reg, col_reg}<16'b0101100101100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101100101100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100101100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101100101100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100101100100) && ({row_reg, col_reg}<16'b0101100101101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100101101000) && ({row_reg, col_reg}<16'b0101100101101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101100101101010) && ({row_reg, col_reg}<16'b0101100101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100101101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100101101101) && ({row_reg, col_reg}<16'b0101100101110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100101110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100101110001) && ({row_reg, col_reg}<16'b0101100101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100101110110) && ({row_reg, col_reg}<16'b0101100101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100101111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101100101111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101100101111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100101111110) && ({row_reg, col_reg}<16'b0101100110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100110000000) && ({row_reg, col_reg}<16'b0101100110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100110000011) && ({row_reg, col_reg}<16'b0101100110101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101100110101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100110101001) && ({row_reg, col_reg}<16'b0101100110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100110101011) && ({row_reg, col_reg}<16'b0101100110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100110110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100110110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100110110010) && ({row_reg, col_reg}<16'b0101100110110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100110110101) && ({row_reg, col_reg}<16'b0101100110111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100110111001) && ({row_reg, col_reg}<16'b0101100110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100110111110) && ({row_reg, col_reg}<16'b0101100111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100111000000) && ({row_reg, col_reg}<16'b0101100111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100111000011) && ({row_reg, col_reg}<16'b0101100111001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100111001101) && ({row_reg, col_reg}<16'b0101100111001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101100111001111) && ({row_reg, col_reg}<16'b0101100111010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100111010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100111010011) && ({row_reg, col_reg}<16'b0101100111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100111011111) && ({row_reg, col_reg}<16'b0101100111100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101100111100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100111100010) && ({row_reg, col_reg}<16'b0101100111100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100111100100) && ({row_reg, col_reg}<16'b0101100111100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100111100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100111100111) && ({row_reg, col_reg}<16'b0101100111110001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0101100111110001) && ({row_reg, col_reg}<16'b0101101000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101101000000000) && ({row_reg, col_reg}<16'b0101101000000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101000000010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0101101000000011) && ({row_reg, col_reg}<16'b0101101000000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101101000000101) && ({row_reg, col_reg}<16'b0101101000000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101101000000111) && ({row_reg, col_reg}<16'b0101101000001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101000001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101101000001011) && ({row_reg, col_reg}<16'b0101101000001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101000001101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0101101000001110) && ({row_reg, col_reg}<16'b0101101000111100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101000111100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0101101000111101) && ({row_reg, col_reg}<16'b0101101000111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101101000111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101001000000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101101001000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101101001000010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101101001000011) && ({row_reg, col_reg}<16'b0101101001000101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101101001000101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101101001000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101101001000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101001001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101001001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101101001001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101001001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101101001001100) && ({row_reg, col_reg}<16'b0101101001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101001001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101001010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101101001010001) && ({row_reg, col_reg}<16'b0101101001010011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101101001010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101101001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101001010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101001010110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101101001010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101001011000) && ({row_reg, col_reg}<16'b0101101001011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101101001011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101001011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101001011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101101001011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101101001011111) && ({row_reg, col_reg}<16'b0101101001100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101001100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101001100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101101001100011) && ({row_reg, col_reg}<16'b0101101001100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101001100101) && ({row_reg, col_reg}<16'b0101101001101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101001101000) && ({row_reg, col_reg}<16'b0101101001101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101101001101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101001101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101001101101) && ({row_reg, col_reg}<16'b0101101001101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101001101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101001110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101001110001) && ({row_reg, col_reg}<16'b0101101001110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101101001110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101001110111) && ({row_reg, col_reg}<16'b0101101001111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101001111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101001111100) && ({row_reg, col_reg}<16'b0101101010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101010000000) && ({row_reg, col_reg}<16'b0101101010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101010000011) && ({row_reg, col_reg}<16'b0101101010101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101101010101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101010101001) && ({row_reg, col_reg}<16'b0101101010101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101010101011) && ({row_reg, col_reg}<16'b0101101010101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101010101111) && ({row_reg, col_reg}<16'b0101101010110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101010110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101010110010) && ({row_reg, col_reg}<16'b0101101010110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101101010110101) && ({row_reg, col_reg}<16'b0101101010111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101010111001) && ({row_reg, col_reg}<16'b0101101010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101010111110) && ({row_reg, col_reg}<16'b0101101011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101011000000) && ({row_reg, col_reg}<16'b0101101011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101101011000011) && ({row_reg, col_reg}<16'b0101101011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101011001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101101011001111) && ({row_reg, col_reg}<16'b0101101011010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101011010011) && ({row_reg, col_reg}<16'b0101101011010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101011010101) && ({row_reg, col_reg}<16'b0101101011011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101011011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101101011011101) && ({row_reg, col_reg}<16'b0101101011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101011011111) && ({row_reg, col_reg}<16'b0101101011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101101011100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101011100010) && ({row_reg, col_reg}<16'b0101101011100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101011100100) && ({row_reg, col_reg}<16'b0101101011100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101011100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101011100111) && ({row_reg, col_reg}<16'b0101101011110001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0101101011110001) && ({row_reg, col_reg}<16'b0101101100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101101100000000) && ({row_reg, col_reg}<16'b0101101100000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101101100000010) && ({row_reg, col_reg}<16'b0101101100000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101101100000101) && ({row_reg, col_reg}<16'b0101101100001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101100001001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0101101100001010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101101100001011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0101101100001100) && ({row_reg, col_reg}<16'b0101101100010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101101100010010) && ({row_reg, col_reg}<16'b0101101100010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0101101100010100) && ({row_reg, col_reg}<16'b0101101100011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101100011000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0101101100011001) && ({row_reg, col_reg}<16'b0101101100100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101101100100000) && ({row_reg, col_reg}<16'b0101101100100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0101101100100010) && ({row_reg, col_reg}<16'b0101101100111100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101100111100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101101100111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101101100111110) && ({row_reg, col_reg}<16'b0101101101000000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101101101000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101101101000001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101101101000010) && ({row_reg, col_reg}<16'b0101101101000101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101101101000101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0101101101000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101101101000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101101001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101101001001) && ({row_reg, col_reg}<16'b0101101101001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101101001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101101101001100) && ({row_reg, col_reg}<16'b0101101101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101101001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101101010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101101101010001) && ({row_reg, col_reg}<16'b0101101101010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101101101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101101010101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101101101010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101101010111) && ({row_reg, col_reg}<16'b0101101101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101101101011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101101011100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101101101011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101101101011110) && ({row_reg, col_reg}<16'b0101101101100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101101100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101101100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101101101100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101101100100) && ({row_reg, col_reg}<16'b0101101101101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101101101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101101101101001) && ({row_reg, col_reg}<16'b0101101101101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101101101101011) && ({row_reg, col_reg}<16'b0101101101101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101101101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101101101101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101101101101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101101110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101101110001) && ({row_reg, col_reg}<16'b0101101101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101101101110110) && ({row_reg, col_reg}<16'b0101101101111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101101101111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101101101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101101101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101110000000) && ({row_reg, col_reg}<16'b0101101110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101110000011) && ({row_reg, col_reg}<16'b0101101110101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101101110101000) && ({row_reg, col_reg}<16'b0101101110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101110101011) && ({row_reg, col_reg}<16'b0101101110101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101110101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101110110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101110110001) && ({row_reg, col_reg}<16'b0101101110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101101110111000) && ({row_reg, col_reg}<16'b0101101110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101110111110) && ({row_reg, col_reg}<16'b0101101111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101111000000) && ({row_reg, col_reg}<16'b0101101111000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101101111000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101111000011) && ({row_reg, col_reg}<16'b0101101111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101111011111) && ({row_reg, col_reg}<16'b0101101111100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101101111100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101111100010) && ({row_reg, col_reg}<16'b0101101111100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101111100100) && ({row_reg, col_reg}<16'b0101101111100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101111100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101111100111) && ({row_reg, col_reg}<16'b0101101111110001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0101101111110001) && ({row_reg, col_reg}<16'b0101110000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101110000000000) && ({row_reg, col_reg}<16'b0101110000000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101110000000010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101110000000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101110000000100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101110000000101) && ({row_reg, col_reg}<16'b0101110000001010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101110000001010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101110000001011) && ({row_reg, col_reg}<16'b0101110000111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101110000111110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0101110000111111) && ({row_reg, col_reg}<16'b0101110001000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101110001000001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101110001000010) && ({row_reg, col_reg}<16'b0101110001000101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101110001000101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101110001000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101110001000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110001001000) && ({row_reg, col_reg}<16'b0101110001001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110001001011) && ({row_reg, col_reg}<16'b0101110001001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110001001101) && ({row_reg, col_reg}<16'b0101110001001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101110001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110001010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101110001010001) && ({row_reg, col_reg}<16'b0101110001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101110001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101110001010101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101110001010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110001010111) && ({row_reg, col_reg}<16'b0101110001011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101110001011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101110001011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101110001011100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101110001011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110001011110) && ({row_reg, col_reg}<16'b0101110001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101110001100010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101110001100011) && ({row_reg, col_reg}<16'b0101110001100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101110001100110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101110001100111) && ({row_reg, col_reg}<16'b0101110001101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101110001101001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101110001101010) && ({row_reg, col_reg}<16'b0101110001101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101110001101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101110001101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110001101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101110001101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110001110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110001110001) && ({row_reg, col_reg}<16'b0101110001110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101110001110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110001110110) && ({row_reg, col_reg}<16'b0101110001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110001111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101110001111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101110001111101) && ({row_reg, col_reg}<16'b0101110010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110010000000) && ({row_reg, col_reg}<16'b0101110010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110010000011) && ({row_reg, col_reg}<16'b0101110010101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101110010101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101110010101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110010101010) && ({row_reg, col_reg}<16'b0101110010101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110010101100) && ({row_reg, col_reg}<16'b0101110010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101110010110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110010110001) && ({row_reg, col_reg}<16'b0101110010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101110010111000) && ({row_reg, col_reg}<16'b0101110010111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110010111010) && ({row_reg, col_reg}<16'b0101110010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110010111110) && ({row_reg, col_reg}<16'b0101110011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110011000000) && ({row_reg, col_reg}<16'b0101110011000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110011000010) && ({row_reg, col_reg}<16'b0101110011000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110011000100) && ({row_reg, col_reg}<16'b0101110011000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110011000110) && ({row_reg, col_reg}<16'b0101110011001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110011001100) && ({row_reg, col_reg}<16'b0101110011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110011011111) && ({row_reg, col_reg}<16'b0101110011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101110011100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110011100010) && ({row_reg, col_reg}<16'b0101110011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110011100111) && ({row_reg, col_reg}<16'b0101110011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110011101111) && ({row_reg, col_reg}<16'b0101110011110001)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0101110011110001) && ({row_reg, col_reg}<16'b0101110100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101110100000000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0101110100000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101110100000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101110100000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101110100000100) && ({row_reg, col_reg}<16'b0101110100000110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101110100000110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101110100000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101110100001000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101110100001001) && ({row_reg, col_reg}<16'b0101110100001100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101110100001100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0101110100001101) && ({row_reg, col_reg}<16'b0101110100010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101110100010000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101110100010001) && ({row_reg, col_reg}<16'b0101110100010100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101110100010100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0101110100010101) && ({row_reg, col_reg}<16'b0101110100011001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101110100011001) && ({row_reg, col_reg}<16'b0101110100100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101110100100011) && ({row_reg, col_reg}<16'b0101110100100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101110100100101) && ({row_reg, col_reg}<16'b0101110100101000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101110100101000) && ({row_reg, col_reg}<16'b0101110100101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101110100101010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101110100101011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101110100101100) && ({row_reg, col_reg}<16'b0101110100110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101110100110101) && ({row_reg, col_reg}<16'b0101110100110111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101110100110111) && ({row_reg, col_reg}<16'b0101110100111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101110100111010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101110100111011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101110100111100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101110100111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101110100111110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0101110100111111) && ({row_reg, col_reg}<16'b0101110101000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101110101000001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101110101000010) && ({row_reg, col_reg}<16'b0101110101000100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101110101000100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0101110101000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101110101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101110101000111) && ({row_reg, col_reg}<16'b0101110101001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101110101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110101001100) && ({row_reg, col_reg}<16'b0101110101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101110101010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101110101010001) && ({row_reg, col_reg}<16'b0101110101010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101110101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101110101010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101110101010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110101010111) && ({row_reg, col_reg}<16'b0101110101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101110101011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110101011100) && ({row_reg, col_reg}<16'b0101110101011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110101011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110101011111) && ({row_reg, col_reg}<16'b0101110101100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101110101100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110101100010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101110101100011) && ({row_reg, col_reg}<16'b0101110101100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110101100110) && ({row_reg, col_reg}<16'b0101110101101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101110101101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110101101010) && ({row_reg, col_reg}<16'b0101110101101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101110101101100) && ({row_reg, col_reg}<16'b0101110101101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110101101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101110101101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110101110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110101110001) && ({row_reg, col_reg}<16'b0101110101110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101110101110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110101110110) && ({row_reg, col_reg}<16'b0101110101111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110101111010) && ({row_reg, col_reg}<16'b0101110101111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110101111101) && ({row_reg, col_reg}<16'b0101110110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110110000011) && ({row_reg, col_reg}<16'b0101110110101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101110110101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101110110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110110101010) && ({row_reg, col_reg}<16'b0101110110101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101110110101101) && ({row_reg, col_reg}<16'b0101110110101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110110101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110110110000) && ({row_reg, col_reg}<16'b0101110110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101110110111000) && ({row_reg, col_reg}<16'b0101110110111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110110111010) && ({row_reg, col_reg}<16'b0101110111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110111000111) && ({row_reg, col_reg}<16'b0101110111001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110111001001) && ({row_reg, col_reg}<16'b0101110111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110111011111) && ({row_reg, col_reg}<16'b0101110111100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101110111100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110111100010) && ({row_reg, col_reg}<16'b0101110111100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110111100111) && ({row_reg, col_reg}<16'b0101110111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110111101111) && ({row_reg, col_reg}<16'b0101110111110001)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0101110111110001) && ({row_reg, col_reg}<16'b0101111000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111000000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101111000000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101111000000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101111000000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101111000000100) && ({row_reg, col_reg}<16'b0101111000000111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101111000000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0101111000001000) && ({row_reg, col_reg}<16'b0101111000001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101111000001101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101111000001110) && ({row_reg, col_reg}<16'b0101111000010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101111000010001) && ({row_reg, col_reg}<16'b0101111000010100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101111000010100) && ({row_reg, col_reg}<16'b0101111000010110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101111000010110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101111000010111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101111000011000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0101111000011001) && ({row_reg, col_reg}<16'b0101111000100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101111000100011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101111000100100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101111000100101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0101111000100110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101111000100111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0101111000101000) && ({row_reg, col_reg}<16'b0101111000101011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101111000101011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0101111000101100) && ({row_reg, col_reg}<16'b0101111000110110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101111000110110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101111000110111) && ({row_reg, col_reg}<16'b0101111000111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101111000111010) && ({row_reg, col_reg}<16'b0101111000111101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101111000111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101111000111110) && ({row_reg, col_reg}<16'b0101111001000000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101111001000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101111001000001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101111001000010) && ({row_reg, col_reg}<16'b0101111001000100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101111001000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101111001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101111001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111001000111) && ({row_reg, col_reg}<16'b0101111001001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101111001001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101111001001100) && ({row_reg, col_reg}<16'b0101111001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101111001010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0101111001010001) && ({row_reg, col_reg}<16'b0101111001010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101111001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101111001010101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101111001010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101111001010111) && ({row_reg, col_reg}<16'b0101111001011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111001011001) && ({row_reg, col_reg}<16'b0101111001011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111001011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101111001011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111001011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101111001011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101111001100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101111001100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101111001100010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101111001100011) && ({row_reg, col_reg}<16'b0101111001100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101111001100110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101111001100111) && ({row_reg, col_reg}<16'b0101111001101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101111001101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101111001101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101111001101011) && ({row_reg, col_reg}<16'b0101111001101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101111001101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101111001101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111001110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111001110001) && ({row_reg, col_reg}<16'b0101111001110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111001110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111001110110) && ({row_reg, col_reg}<16'b0101111001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111001111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111001111100) && ({row_reg, col_reg}<16'b0101111001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111001111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111010000001) && ({row_reg, col_reg}<16'b0101111010000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111010000011) && ({row_reg, col_reg}<16'b0101111010101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111010101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111010101010) && ({row_reg, col_reg}<16'b0101111010101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111010101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101111010101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111010110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111010110001) && ({row_reg, col_reg}<16'b0101111010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101111010111000) && ({row_reg, col_reg}<16'b0101111011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111011000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101111011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101111011000010) && ({row_reg, col_reg}<16'b0101111011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111011001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101111011001001) && ({row_reg, col_reg}<16'b0101111011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111011011111) && ({row_reg, col_reg}<16'b0101111011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111011100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111011100010) && ({row_reg, col_reg}<16'b0101111011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101111011100111) && ({row_reg, col_reg}<16'b0101111011101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111011101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111011101010) && ({row_reg, col_reg}<16'b0101111011110001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0101111011110001) && ({row_reg, col_reg}<16'b0101111100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111100000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101111100000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101111100000010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101111100000011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101111100000100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0101111100000101) && ({row_reg, col_reg}<16'b0101111100001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101111100001101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0101111100001110) && ({row_reg, col_reg}<16'b0101111100010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101111100010010) && ({row_reg, col_reg}<16'b0101111100010100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101111100010100) && ({row_reg, col_reg}<16'b0101111100010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101111100010110) && ({row_reg, col_reg}<16'b0101111100011001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101111100011001) && ({row_reg, col_reg}<16'b0101111100100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101111100100100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101111100100101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0101111100100110) && ({row_reg, col_reg}<16'b0101111100101011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101111100101011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0101111100101100) && ({row_reg, col_reg}<16'b0101111100110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101111100110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101111100110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101111100110111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101111100111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101111100111001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101111100111010) && ({row_reg, col_reg}<16'b0101111100111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101111100111110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101111100111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101111101000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101111101000001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101111101000010)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0101111101000011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101111101000100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101111101000101) && ({row_reg, col_reg}<16'b0101111101000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111101000111) && ({row_reg, col_reg}<16'b0101111101001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101111101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111101001100) && ({row_reg, col_reg}<16'b0101111101001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101111101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101111101010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101111101010001) && ({row_reg, col_reg}<16'b0101111101010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101111101010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101111101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101111101010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111101010110) && ({row_reg, col_reg}<16'b0101111101011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101111101011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111101011001) && ({row_reg, col_reg}<16'b0101111101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111101011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101111101011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111101011101) && ({row_reg, col_reg}<16'b0101111101011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101111101011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101111101100000)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}==16'b0101111101100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101111101100010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101111101100011) && ({row_reg, col_reg}<16'b0101111101100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101111101100110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101111101100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101111101101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101111101101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111101101010) && ({row_reg, col_reg}<16'b0101111101101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101111101101100) && ({row_reg, col_reg}<16'b0101111101101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101111101101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101111101101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111101110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111101110001) && ({row_reg, col_reg}<16'b0101111101110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111101110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111101110110) && ({row_reg, col_reg}<16'b0101111101111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111101111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101111101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111101111100) && ({row_reg, col_reg}<16'b0101111101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111101111110) && ({row_reg, col_reg}<16'b0101111110000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101111110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111110000011) && ({row_reg, col_reg}<16'b0101111110101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111110101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101111110101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111110110000) && ({row_reg, col_reg}<16'b0101111110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101111110111000) && ({row_reg, col_reg}<16'b0101111111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111111000000) && ({row_reg, col_reg}<16'b0101111111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101111111000011) && ({row_reg, col_reg}<16'b0101111111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111111001000) && ({row_reg, col_reg}<16'b0101111111001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101111111001010) && ({row_reg, col_reg}<16'b0101111111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111111011111) && ({row_reg, col_reg}<16'b0101111111100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111111100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111111100010) && ({row_reg, col_reg}<16'b0101111111100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101111111100111) && ({row_reg, col_reg}<16'b0101111111110001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0101111111110001) && ({row_reg, col_reg}<16'b0110000000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110000000000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110000000000001) && ({row_reg, col_reg}<16'b0110000000000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110000000000110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110000000000111) && ({row_reg, col_reg}<16'b0110000000001011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110000000001011) && ({row_reg, col_reg}<16'b0110000000001111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110000000001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110000000010000) && ({row_reg, col_reg}<16'b0110000000010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000000010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110000000010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110000000010100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110000000010101) && ({row_reg, col_reg}<16'b0110000000011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110000000011010) && ({row_reg, col_reg}<16'b0110000000011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110000000011100) && ({row_reg, col_reg}<16'b0110000000011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110000000011110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110000000011111) && ({row_reg, col_reg}<16'b0110000000100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110000000100001) && ({row_reg, col_reg}<16'b0110000000100110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110000000100110) && ({row_reg, col_reg}<16'b0110000000101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110000000101010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110000000101011) && ({row_reg, col_reg}<16'b0110000000101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110000000101111) && ({row_reg, col_reg}<16'b0110000000111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110000000111010) && ({row_reg, col_reg}<16'b0110000000111100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110000000111100) && ({row_reg, col_reg}<16'b0110000001000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110000001000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110000001000001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110000001000010)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0110000001000011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110000001000100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110000001000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110000001000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0110000001000111) && ({row_reg, col_reg}<16'b0110000001001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110000001001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110000001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110000001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000001001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110000001001110) && ({row_reg, col_reg}<16'b0110000001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000001010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0110000001010001) && ({row_reg, col_reg}<16'b0110000001010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110000001010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110000001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000001010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110000001010110) && ({row_reg, col_reg}<16'b0110000001011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110000001011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000001011010) && ({row_reg, col_reg}<16'b0110000001011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000001011100) && ({row_reg, col_reg}<16'b0110000001011110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110000001011110) && ({row_reg, col_reg}<16'b0110000001100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110000001100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000001100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110000001100010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110000001100011) && ({row_reg, col_reg}<16'b0110000001100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000001100110) && ({row_reg, col_reg}<16'b0110000001101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110000001101000) && ({row_reg, col_reg}<16'b0110000001101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110000001101010) && ({row_reg, col_reg}<16'b0110000001101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110000001101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110000001101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000001110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000001110001) && ({row_reg, col_reg}<16'b0110000001110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110000001110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000001110110) && ({row_reg, col_reg}<16'b0110000001111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000001111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000001111011) && ({row_reg, col_reg}<16'b0110000001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000001111110) && ({row_reg, col_reg}<16'b0110000010000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110000010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110000010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000010000011) && ({row_reg, col_reg}<16'b0110000010101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110000010101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110000010101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000010110000) && ({row_reg, col_reg}<16'b0110000010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110000010111000) && ({row_reg, col_reg}<16'b0110000010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000010111110) && ({row_reg, col_reg}<16'b0110000011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000011000000) && ({row_reg, col_reg}<16'b0110000011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110000011000011) && ({row_reg, col_reg}<16'b0110000011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000011001000) && ({row_reg, col_reg}<16'b0110000011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000011001011) && ({row_reg, col_reg}<16'b0110000011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000011011111) && ({row_reg, col_reg}<16'b0110000011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110000011100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000011100010) && ({row_reg, col_reg}<16'b0110000011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000011100111) && ({row_reg, col_reg}<16'b0110000011110001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0110000011110001) && ({row_reg, col_reg}<16'b0110000100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110000100000000) && ({row_reg, col_reg}<16'b0110000100000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110000100000011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110000100000100) && ({row_reg, col_reg}<16'b0110000100000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000100000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110000100000111) && ({row_reg, col_reg}<16'b0110000100001011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110000100001011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110000100001100) && ({row_reg, col_reg}<16'b0110000100001111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110000100001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110000100010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000100010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110000100010010) && ({row_reg, col_reg}<16'b0110000100011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000100011001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110000100011010) && ({row_reg, col_reg}<16'b0110000100100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110000100100011) && ({row_reg, col_reg}<16'b0110000100100110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110000100100110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110000100100111) && ({row_reg, col_reg}<16'b0110000100101001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110000100101001) && ({row_reg, col_reg}<16'b0110000100101101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110000100101101) && ({row_reg, col_reg}<16'b0110000100110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110000100110000) && ({row_reg, col_reg}<16'b0110000100110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110000100110111) && ({row_reg, col_reg}<16'b0110000100111001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110000100111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000100111010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110000100111011) && ({row_reg, col_reg}<16'b0110000100111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110000100111110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110000100111111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110000101000000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0110000101000001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110000101000010)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==16'b0110000101000011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110000101000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110000101000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110000101000110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0110000101000111) && ({row_reg, col_reg}<16'b0110000101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000101001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110000101001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000101001100)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0110000101001101) && ({row_reg, col_reg}<16'b0110000101001111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110000101001111) && ({row_reg, col_reg}<16'b0110000101010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110000101010010)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0110000101010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110000101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000101010101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110000101010110) && ({row_reg, col_reg}<16'b0110000101011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110000101011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110000101011100) && ({row_reg, col_reg}<16'b0110000101100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110000101100000) && ({row_reg, col_reg}<16'b0110000101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110000101100010) && ({row_reg, col_reg}<16'b0110000101100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110000101100100) && ({row_reg, col_reg}<16'b0110000101100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000101100110) && ({row_reg, col_reg}<16'b0110000101101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110000101101000) && ({row_reg, col_reg}<16'b0110000101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110000101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110000101101011) && ({row_reg, col_reg}<16'b0110000101101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110000101101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110000101101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110000101101111) && ({row_reg, col_reg}<16'b0110000101110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000101110001) && ({row_reg, col_reg}<16'b0110000101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110000101110110) && ({row_reg, col_reg}<16'b0110000101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000101111011) && ({row_reg, col_reg}<16'b0110000101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110000101111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110000110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110000110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000110000011) && ({row_reg, col_reg}<16'b0110000110100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110000110100111) && ({row_reg, col_reg}<16'b0110000110101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000110101010) && ({row_reg, col_reg}<16'b0110000110101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110000110101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110000110101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000110110000) && ({row_reg, col_reg}<16'b0110000110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110000110111000) && ({row_reg, col_reg}<16'b0110000110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000110111110) && ({row_reg, col_reg}<16'b0110000111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000111000000) && ({row_reg, col_reg}<16'b0110000111000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110000111000010)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==16'b0110000111000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000111000100) && ({row_reg, col_reg}<16'b0110000111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000111001000) && ({row_reg, col_reg}<16'b0110000111001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000111001100) && ({row_reg, col_reg}<16'b0110000111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000111011111) && ({row_reg, col_reg}<16'b0110000111100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000111100010) && ({row_reg, col_reg}<16'b0110000111110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000111110000)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0110000111110001) && ({row_reg, col_reg}<16'b0110001000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110001000000000) && ({row_reg, col_reg}<16'b0110001000000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001000000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110001000000100) && ({row_reg, col_reg}<16'b0110001000000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001000000110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0110001000000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001000001000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110001000001001) && ({row_reg, col_reg}<16'b0110001000001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001000001110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110001000001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001000010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001000010001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0110001000010010) && ({row_reg, col_reg}<16'b0110001000011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001000011011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110001000011100) && ({row_reg, col_reg}<16'b0110001000011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001000011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110001000011111) && ({row_reg, col_reg}<16'b0110001000100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110001000100010) && ({row_reg, col_reg}<16'b0110001000101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001000101111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110001000110000) && ({row_reg, col_reg}<16'b0110001000110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110001000110110) && ({row_reg, col_reg}<16'b0110001000111001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110001000111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001000111010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110001000111011) && ({row_reg, col_reg}<16'b0110001000111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001000111101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110001000111110)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0110001000111111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0110001001000000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0110001001000001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110001001000010)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0110001001000011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110001001000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110001001000101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110001001000110) && ({row_reg, col_reg}<16'b0110001001001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001001001011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110001001001100) && ({row_reg, col_reg}<16'b0110001001010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110001001010000) && ({row_reg, col_reg}<16'b0110001001010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110001001010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001001010101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110001001010110) && ({row_reg, col_reg}<16'b0110001001011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110001001011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001001011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001001011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110001001011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110001001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001001100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001001100001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0110001001100010) && ({row_reg, col_reg}<16'b0110001001100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110001001100100) && ({row_reg, col_reg}<16'b0110001001100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110001001100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110001001101000) && ({row_reg, col_reg}<16'b0110001001101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001001101010) && ({row_reg, col_reg}<16'b0110001001101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110001001101100) && ({row_reg, col_reg}<16'b0110001001110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110001001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001001110001) && ({row_reg, col_reg}<16'b0110001001110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110001001110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001001110111) && ({row_reg, col_reg}<16'b0110001001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001001111011) && ({row_reg, col_reg}<16'b0110001001111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001001111101) && ({row_reg, col_reg}<16'b0110001001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001010000000) && ({row_reg, col_reg}<16'b0110001010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001010000011) && ({row_reg, col_reg}<16'b0110001010100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110001010100100) && ({row_reg, col_reg}<16'b0110001010101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001010101000) && ({row_reg, col_reg}<16'b0110001010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001010101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001010101011) && ({row_reg, col_reg}<16'b0110001010101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110001010101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001010101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110001010110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001010110001) && ({row_reg, col_reg}<16'b0110001010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110001010111000) && ({row_reg, col_reg}<16'b0110001010111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001010111010) && ({row_reg, col_reg}<16'b0110001010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001010111110) && ({row_reg, col_reg}<16'b0110001011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001011000000) && ({row_reg, col_reg}<16'b0110001011000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001011000010) && ({row_reg, col_reg}<16'b0110001011000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001011000100) && ({row_reg, col_reg}<16'b0110001011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001011001000) && ({row_reg, col_reg}<16'b0110001011001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001011001101) && ({row_reg, col_reg}<16'b0110001011010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001011010110) && ({row_reg, col_reg}<16'b0110001011011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001011011000) && ({row_reg, col_reg}<16'b0110001011011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001011011100) && ({row_reg, col_reg}<16'b0110001011011110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110001011011110) && ({row_reg, col_reg}<16'b0110001011100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001011100000) && ({row_reg, col_reg}<16'b0110001011100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001011100010) && ({row_reg, col_reg}<16'b0110001011110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001011110000)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0110001011110001) && ({row_reg, col_reg}<16'b0110001100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110001100000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001100000001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110001100000010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001100000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001100000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110001100000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110001100000111) && ({row_reg, col_reg}<16'b0110001100001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001100001001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110001100001010) && ({row_reg, col_reg}<16'b0110001100001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110001100001101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110001100001110) && ({row_reg, col_reg}<16'b0110001100010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001100010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001100010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110001100010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110001100010011) && ({row_reg, col_reg}<16'b0110001100010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001100010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110001100010111) && ({row_reg, col_reg}<16'b0110001100011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001100011001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110001100011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001100011011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110001100011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001100011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110001100011110) && ({row_reg, col_reg}<16'b0110001100100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110001100100101) && ({row_reg, col_reg}<16'b0110001100101001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110001100101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110001100101010) && ({row_reg, col_reg}<16'b0110001100101110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110001100101110) && ({row_reg, col_reg}<16'b0110001100110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110001100110000) && ({row_reg, col_reg}<16'b0110001100110011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110001100110011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110001100110100) && ({row_reg, col_reg}<16'b0110001100111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001100111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110001100111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110001100111101) && ({row_reg, col_reg}<16'b0110001100111111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110001100111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001101000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110001101000001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110001101000010)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0110001101000011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110001101000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110001101000101) && ({row_reg, col_reg}<16'b0110001101001001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110001101001001) && ({row_reg, col_reg}<16'b0110001101001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001101001111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110001101010000) && ({row_reg, col_reg}<16'b0110001101010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001101010010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0110001101010011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110001101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001101010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001101010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110001101010111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110001101011000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110001101011001) && ({row_reg, col_reg}<16'b0110001101011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001101011011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110001101011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001101011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110001101011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110001101011111) && ({row_reg, col_reg}<16'b0110001101100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001101100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001101100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110001101100011) && ({row_reg, col_reg}<16'b0110001101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001101101011) && ({row_reg, col_reg}<16'b0110001101101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001101101101) && ({row_reg, col_reg}<16'b0110001101101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110001101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110001101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001101110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001101110010) && ({row_reg, col_reg}<16'b0110001101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110001101110110) && ({row_reg, col_reg}<16'b0110001110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001110000011) && ({row_reg, col_reg}<16'b0110001110100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110001110100100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001110100101) && ({row_reg, col_reg}<16'b0110001110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001110101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110001110101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110001110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001110101110) && ({row_reg, col_reg}<16'b0110001110110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001110110001) && ({row_reg, col_reg}<16'b0110001110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110001110111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001110111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001110111010) && ({row_reg, col_reg}<16'b0110001110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001110111110) && ({row_reg, col_reg}<16'b0110001111000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001111000001) && ({row_reg, col_reg}<16'b0110001111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001111000111) && ({row_reg, col_reg}<16'b0110001111001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001111001101) && ({row_reg, col_reg}<16'b0110001111011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001111011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001111011010) && ({row_reg, col_reg}<16'b0110001111011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001111011100) && ({row_reg, col_reg}<16'b0110001111011110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110001111011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001111011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110001111100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110001111100001) && ({row_reg, col_reg}<16'b0110001111110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001111110000)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0110001111110001) && ({row_reg, col_reg}<16'b0110010000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110010000000000) && ({row_reg, col_reg}<16'b0110010000000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110010000000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110010000000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010000000101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110010000000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110010000000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110010000001000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110010000001001) && ({row_reg, col_reg}<16'b0110010000001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110010000001110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110010000001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110010000010000) && ({row_reg, col_reg}<16'b0110010000010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110010000010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110010000010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110010000010100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110010000010101) && ({row_reg, col_reg}<16'b0110010000011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110010000011000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110010000011001) && ({row_reg, col_reg}<16'b0110010000011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110010000011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110010000011111) && ({row_reg, col_reg}<16'b0110010000100001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110010000100001)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0110010000100010) && ({row_reg, col_reg}<16'b0110010000100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110010000100101) && ({row_reg, col_reg}<16'b0110010000101001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110010000101001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110010000101010) && ({row_reg, col_reg}<16'b0110010000101111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110010000101111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110010000110000) && ({row_reg, col_reg}<16'b0110010000110100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110010000110100) && ({row_reg, col_reg}<16'b0110010000110110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110010000110110) && ({row_reg, col_reg}<16'b0110010000111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110010000111010) && ({row_reg, col_reg}<16'b0110010000111100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110010000111100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110010000111101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0110010000111110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110010000111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110010001000000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110010001000001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0110010001000010) && ({row_reg, col_reg}<16'b0110010001000100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0110010001000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110010001000101) && ({row_reg, col_reg}<16'b0110010001001000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110010001001000) && ({row_reg, col_reg}<16'b0110010001001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110010001001101) && ({row_reg, col_reg}<16'b0110010001010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110010001010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110010001010111) && ({row_reg, col_reg}<16'b0110010001011001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110010001011001) && ({row_reg, col_reg}<16'b0110010001011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010001011011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110010001011100) && ({row_reg, col_reg}<16'b0110010001011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110010001011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110010001011111) && ({row_reg, col_reg}<16'b0110010001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110010001100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110010001100011) && ({row_reg, col_reg}<16'b0110010001101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110010001101011) && ({row_reg, col_reg}<16'b0110010001101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010001101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110010001101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110010001101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010001110001) && ({row_reg, col_reg}<16'b0110010001110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110010001110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110010001110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010001110111) && ({row_reg, col_reg}<16'b0110010010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010010000010) && ({row_reg, col_reg}<16'b0110010010100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110010010100100) && ({row_reg, col_reg}<16'b0110010010100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010010100111) && ({row_reg, col_reg}<16'b0110010010101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010010101001) && ({row_reg, col_reg}<16'b0110010010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010010101101) && ({row_reg, col_reg}<16'b0110010010110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110010010110001) && ({row_reg, col_reg}<16'b0110010010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110010010111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010010111001) && ({row_reg, col_reg}<16'b0110010010111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010010111111) && ({row_reg, col_reg}<16'b0110010011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010011000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010011000010) && ({row_reg, col_reg}<16'b0110010011000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010011000110) && ({row_reg, col_reg}<16'b0110010011001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110010011001101) && ({row_reg, col_reg}<16'b0110010011010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010011010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010011010101) && ({row_reg, col_reg}<16'b0110010011011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010011011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110010011011010) && ({row_reg, col_reg}<16'b0110010011011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010011011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110010011011101) && ({row_reg, col_reg}<16'b0110010011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010011011111) && ({row_reg, col_reg}<16'b0110010011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110010011100001) && ({row_reg, col_reg}<16'b0110010011110001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0110010011110001) && ({row_reg, col_reg}<16'b0110010100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110010100000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110010100000001) && ({row_reg, col_reg}<16'b0110010100000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110010100000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110010100000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010100000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110010100000110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110010100000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110010100001000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110010100001001) && ({row_reg, col_reg}<16'b0110010100001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110010100001011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110010100001100) && ({row_reg, col_reg}<16'b0110010100001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110010100001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110010100001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110010100010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110010100010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110010100010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110010100010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110010100010100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110010100010101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110010100010110) && ({row_reg, col_reg}<16'b0110010100011101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110010100011101) && ({row_reg, col_reg}<16'b0110010100100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110010100100011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110010100100100) && ({row_reg, col_reg}<16'b0110010100110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110010100110010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110010100110011) && ({row_reg, col_reg}<16'b0110010100110110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110010100110110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110010100110111) && ({row_reg, col_reg}<16'b0110010100111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110010100111001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110010100111010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110010100111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110010100111100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110010100111101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110010100111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110010100111111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110010101000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110010101000001) && ({row_reg, col_reg}<16'b0110010101000100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110010101000100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110010101000101) && ({row_reg, col_reg}<16'b0110010101001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110010101001001) && ({row_reg, col_reg}<16'b0110010101001011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110010101001011) && ({row_reg, col_reg}<16'b0110010101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110010101010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110010101010101) && ({row_reg, col_reg}<16'b0110010101010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110010101010111) && ({row_reg, col_reg}<16'b0110010101011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110010101011100) && ({row_reg, col_reg}<16'b0110010101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110010101011110) && ({row_reg, col_reg}<16'b0110010101100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110010101100000) && ({row_reg, col_reg}<16'b0110010101100010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110010101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110010101100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110010101100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010101100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110010101100110) && ({row_reg, col_reg}<16'b0110010101101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110010101101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110010101101001) && ({row_reg, col_reg}<16'b0110010101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110010101101011) && ({row_reg, col_reg}<16'b0110010101101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010101101101) && ({row_reg, col_reg}<16'b0110010101110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110010101110000) && ({row_reg, col_reg}<16'b0110010101110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010101110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110010101110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110010101110110) && ({row_reg, col_reg}<16'b0110010101111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010101111000) && ({row_reg, col_reg}<16'b0110010101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010101111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010101111100) && ({row_reg, col_reg}<16'b0110010110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010110000010) && ({row_reg, col_reg}<16'b0110010110100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110010110100100) && ({row_reg, col_reg}<16'b0110010110100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110010110100111) && ({row_reg, col_reg}<16'b0110010110101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010110101011) && ({row_reg, col_reg}<16'b0110010110110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110010110110001) && ({row_reg, col_reg}<16'b0110010110110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110010110110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010110110101) && ({row_reg, col_reg}<16'b0110010110110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110010110110111) && ({row_reg, col_reg}<16'b0110010110111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010110111001) && ({row_reg, col_reg}<16'b0110010110111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010110111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010110111101) && ({row_reg, col_reg}<16'b0110010110111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010110111111) && ({row_reg, col_reg}<16'b0110010111000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010111000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010111000010) && ({row_reg, col_reg}<16'b0110010111000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010111000110) && ({row_reg, col_reg}<16'b0110010111001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110010111001000) && ({row_reg, col_reg}<16'b0110010111001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010111001010) && ({row_reg, col_reg}<16'b0110010111001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110010111001101) && ({row_reg, col_reg}<16'b0110010111010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010111010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010111010001) && ({row_reg, col_reg}<16'b0110010111010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010111010011) && ({row_reg, col_reg}<16'b0110010111010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010111010101) && ({row_reg, col_reg}<16'b0110010111011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010111011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110010111011010) && ({row_reg, col_reg}<16'b0110010111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010111011111) && ({row_reg, col_reg}<16'b0110010111100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110010111100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010111100010) && ({row_reg, col_reg}<16'b0110010111100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010111100100) && ({row_reg, col_reg}<16'b0110010111100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110010111100111) && ({row_reg, col_reg}<16'b0110010111101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010111101110) && ({row_reg, col_reg}<16'b0110010111110001)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0110010111110001) && ({row_reg, col_reg}<16'b0110011000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110011000000000) && ({row_reg, col_reg}<16'b0110011000000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110011000000010) && ({row_reg, col_reg}<16'b0110011000000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110011000000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110011000000110) && ({row_reg, col_reg}<16'b0110011000001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011000001110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110011000001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110011000010000) && ({row_reg, col_reg}<16'b0110011000010010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0110011000010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011000010011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110011000010100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110011000010101) && ({row_reg, col_reg}<16'b0110011000011000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110011000011000) && ({row_reg, col_reg}<16'b0110011000011010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110011000011010) && ({row_reg, col_reg}<16'b0110011000011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110011000011100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110011000011101) && ({row_reg, col_reg}<16'b0110011000100000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110011000100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011000100001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110011000100010) && ({row_reg, col_reg}<16'b0110011000100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110011000100101) && ({row_reg, col_reg}<16'b0110011000101000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110011000101000) && ({row_reg, col_reg}<16'b0110011000101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110011000101010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110011000101011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110011000101100) && ({row_reg, col_reg}<16'b0110011000110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110011000110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110011000110001) && ({row_reg, col_reg}<16'b0110011000110111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110011000110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110011000111000) && ({row_reg, col_reg}<16'b0110011000111010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110011000111010) && ({row_reg, col_reg}<16'b0110011000111100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110011000111100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110011000111101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110011000111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011000111111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110011001000000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0110011001000001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110011001000010) && ({row_reg, col_reg}<16'b0110011001000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011001000100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110011001000101) && ({row_reg, col_reg}<16'b0110011001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110011001010100) && ({row_reg, col_reg}<16'b0110011001010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110011001010110) && ({row_reg, col_reg}<16'b0110011001011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110011001011001) && ({row_reg, col_reg}<16'b0110011001011011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0110011001011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110011001011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110011001011101) && ({row_reg, col_reg}<16'b0110011001011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110011001011111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110011001100000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110011001100001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0110011001100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110011001100011) && ({row_reg, col_reg}<16'b0110011001100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110011001100101) && ({row_reg, col_reg}<16'b0110011001101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110011001101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110011001101001) && ({row_reg, col_reg}<16'b0110011001101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110011001101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110011001101101) && ({row_reg, col_reg}<16'b0110011001110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110011001110000) && ({row_reg, col_reg}<16'b0110011001110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011001110011) && ({row_reg, col_reg}<16'b0110011001111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011001111000) && ({row_reg, col_reg}<16'b0110011001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011001111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110011001111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011001111101) && ({row_reg, col_reg}<16'b0110011010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011010000011) && ({row_reg, col_reg}<16'b0110011010100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110011010100100) && ({row_reg, col_reg}<16'b0110011010100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110011010100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011010100111) && ({row_reg, col_reg}<16'b0110011010101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110011010101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110011010101011) && ({row_reg, col_reg}<16'b0110011010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110011010110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011010110001) && ({row_reg, col_reg}<16'b0110011010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110011010111000) && ({row_reg, col_reg}<16'b0110011010111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011010111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011010111101) && ({row_reg, col_reg}<16'b0110011010111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011010111111) && ({row_reg, col_reg}<16'b0110011011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110011011000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011011000010) && ({row_reg, col_reg}<16'b0110011011000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011011000110) && ({row_reg, col_reg}<16'b0110011011001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011011001000) && ({row_reg, col_reg}<16'b0110011011001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011011001011) && ({row_reg, col_reg}<16'b0110011011001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011011001101) && ({row_reg, col_reg}<16'b0110011011010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011011010000) && ({row_reg, col_reg}<16'b0110011011010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011011010010) && ({row_reg, col_reg}<16'b0110011011010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011011010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011011010101) && ({row_reg, col_reg}<16'b0110011011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011011011111) && ({row_reg, col_reg}<16'b0110011011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110011011100001) && ({row_reg, col_reg}<16'b0110011011100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011011100100) && ({row_reg, col_reg}<16'b0110011011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011011100111) && ({row_reg, col_reg}<16'b0110011011101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011011101110) && ({row_reg, col_reg}<16'b0110011011110001)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0110011011110001) && ({row_reg, col_reg}<16'b0110011100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110011100000000) && ({row_reg, col_reg}<16'b0110011100000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110011100000010) && ({row_reg, col_reg}<16'b0110011100000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110011100000100) && ({row_reg, col_reg}<16'b0110011100000110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110011100000110)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0110011100000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110011100001000) && ({row_reg, col_reg}<16'b0110011100001010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110011100001010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110011100001011) && ({row_reg, col_reg}<16'b0110011100001111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110011100001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110011100010000) && ({row_reg, col_reg}<16'b0110011100010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110011100010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011100010011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110011100010100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110011100010101) && ({row_reg, col_reg}<16'b0110011100011000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110011100011000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110011100011001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110011100011010) && ({row_reg, col_reg}<16'b0110011100011101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110011100011101) && ({row_reg, col_reg}<16'b0110011100100001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110011100100001) && ({row_reg, col_reg}<16'b0110011100100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110011100100101) && ({row_reg, col_reg}<16'b0110011100101000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110011100101000) && ({row_reg, col_reg}<16'b0110011100101011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110011100101011) && ({row_reg, col_reg}<16'b0110011100110010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110011100110010) && ({row_reg, col_reg}<16'b0110011100110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011100110111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110011100111000) && ({row_reg, col_reg}<16'b0110011100111011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110011100111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110011100111100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110011100111101) && ({row_reg, col_reg}<16'b0110011100111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011100111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110011101000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110011101000001) && ({row_reg, col_reg}<16'b0110011101000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110011101000011) && ({row_reg, col_reg}<16'b0110011101010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110011101010001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110011101010010) && ({row_reg, col_reg}<16'b0110011101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110011101010100) && ({row_reg, col_reg}<16'b0110011101010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110011101010110) && ({row_reg, col_reg}<16'b0110011101011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110011101011000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110011101011001) && ({row_reg, col_reg}<16'b0110011101011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110011101011111) && ({row_reg, col_reg}<16'b0110011101100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110011101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110011101100011) && ({row_reg, col_reg}<16'b0110011101100110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110011101100110) && ({row_reg, col_reg}<16'b0110011101101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110011101101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110011101101001) && ({row_reg, col_reg}<16'b0110011101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011101101100) && ({row_reg, col_reg}<16'b0110011101101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110011101101110) && ({row_reg, col_reg}<16'b0110011101110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110011101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011101110001) && ({row_reg, col_reg}<16'b0110011101111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011101111000) && ({row_reg, col_reg}<16'b0110011101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011101111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011101111100) && ({row_reg, col_reg}<16'b0110011101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011110000000) && ({row_reg, col_reg}<16'b0110011110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011110000011) && ({row_reg, col_reg}<16'b0110011110100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110011110100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011110100100) && ({row_reg, col_reg}<16'b0110011110100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110011110100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011110100111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011110101000) && ({row_reg, col_reg}<16'b0110011110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011110101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110011110101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110011110101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011110101101) && ({row_reg, col_reg}<16'b0110011110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011110110000) && ({row_reg, col_reg}<16'b0110011110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110011110111000) && ({row_reg, col_reg}<16'b0110011110111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011110111010) && ({row_reg, col_reg}<16'b0110011110111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011110111111) && ({row_reg, col_reg}<16'b0110011111000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110011111000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011111000010) && ({row_reg, col_reg}<16'b0110011111000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011111000110) && ({row_reg, col_reg}<16'b0110011111001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011111001000) && ({row_reg, col_reg}<16'b0110011111001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011111001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011111001101) && ({row_reg, col_reg}<16'b0110011111010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011111010011) && ({row_reg, col_reg}<16'b0110011111010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011111010110) && ({row_reg, col_reg}<16'b0110011111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011111011111) && ({row_reg, col_reg}<16'b0110011111100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110011111100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011111100010) && ({row_reg, col_reg}<16'b0110011111100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011111100111) && ({row_reg, col_reg}<16'b0110011111101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011111101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110011111101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011111101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110011111110000)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0110011111110001) && ({row_reg, col_reg}<16'b0110100000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110100000000000) && ({row_reg, col_reg}<16'b0110100000000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110100000000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110100000000110) && ({row_reg, col_reg}<16'b0110100000001000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110100000001000) && ({row_reg, col_reg}<16'b0110100000001101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110100000001101) && ({row_reg, col_reg}<16'b0110100000001111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110100000001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110100000010000) && ({row_reg, col_reg}<16'b0110100000010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110100000010010) && ({row_reg, col_reg}<16'b0110100000010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110100000010101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110100000010110) && ({row_reg, col_reg}<16'b0110100000011000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110100000011000) && ({row_reg, col_reg}<16'b0110100000011011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110100000011011) && ({row_reg, col_reg}<16'b0110100000011110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110100000011110) && ({row_reg, col_reg}<16'b0110100000100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110100000100001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110100000100010) && ({row_reg, col_reg}<16'b0110100000100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110100000100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110100000100110) && ({row_reg, col_reg}<16'b0110100000101000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110100000101000) && ({row_reg, col_reg}<16'b0110100000101011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110100000101011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110100000101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110100000101101) && ({row_reg, col_reg}<16'b0110100000101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110100000101111) && ({row_reg, col_reg}<16'b0110100000110001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110100000110001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110100000110010) && ({row_reg, col_reg}<16'b0110100000111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110100000111101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110100000111110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110100000111111) && ({row_reg, col_reg}<16'b0110100001000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110100001000001) && ({row_reg, col_reg}<16'b0110100001000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110100001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110100001000110) && ({row_reg, col_reg}<16'b0110100001001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110100001001000) && ({row_reg, col_reg}<16'b0110100001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110100001001100) && ({row_reg, col_reg}<16'b0110100001001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110100001001110) && ({row_reg, col_reg}<16'b0110100001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110100001010000) && ({row_reg, col_reg}<16'b0110100001010111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110100001010111) && ({row_reg, col_reg}<16'b0110100001011001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110100001011001) && ({row_reg, col_reg}<16'b0110100001011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110100001011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110100001011110) && ({row_reg, col_reg}<16'b0110100001100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110100001100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110100001100001) && ({row_reg, col_reg}<16'b0110100001100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110100001100011) && ({row_reg, col_reg}<16'b0110100001100110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110100001100110) && ({row_reg, col_reg}<16'b0110100001101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110100001101000) && ({row_reg, col_reg}<16'b0110100001101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100001101101) && ({row_reg, col_reg}<16'b0110100001101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110100001101111) && ({row_reg, col_reg}<16'b0110100001110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100001110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100001110010) && ({row_reg, col_reg}<16'b0110100001110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110100001110100) && ({row_reg, col_reg}<16'b0110100001111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100001111000) && ({row_reg, col_reg}<16'b0110100001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100001111100) && ({row_reg, col_reg}<16'b0110100001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100001111110) && ({row_reg, col_reg}<16'b0110100010000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110100010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110100010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100010000011) && ({row_reg, col_reg}<16'b0110100010100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110100010100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100010100100) && ({row_reg, col_reg}<16'b0110100010100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100010100111) && ({row_reg, col_reg}<16'b0110100010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100010101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100010101011) && ({row_reg, col_reg}<16'b0110100010101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110100010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100010101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110100010101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100010110000) && ({row_reg, col_reg}<16'b0110100010110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110100010110111) && ({row_reg, col_reg}<16'b0110100010111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100010111010) && ({row_reg, col_reg}<16'b0110100010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100010111110) && ({row_reg, col_reg}<16'b0110100011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100011000001) && ({row_reg, col_reg}<16'b0110100011000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100011000011) && ({row_reg, col_reg}<16'b0110100011010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100011010011) && ({row_reg, col_reg}<16'b0110100011010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100011010111) && ({row_reg, col_reg}<16'b0110100011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100011011111) && ({row_reg, col_reg}<16'b0110100011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110100011100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100011100010) && ({row_reg, col_reg}<16'b0110100011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100011100111) && ({row_reg, col_reg}<16'b0110100011101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100011101100) && ({row_reg, col_reg}<16'b0110100011101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110100011101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100011101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110100011110000)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0110100011110001) && ({row_reg, col_reg}<16'b0110100100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110100100000000) && ({row_reg, col_reg}<16'b0110100100000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110100100000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110100100000110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110100100000111) && ({row_reg, col_reg}<16'b0110100100001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110100100001110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110100100001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110100100010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110100100010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110100100010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110100100010011) && ({row_reg, col_reg}<16'b0110100100010101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110100100010101) && ({row_reg, col_reg}<16'b0110100100011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110100100011011) && ({row_reg, col_reg}<16'b0110100100011110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110100100011110) && ({row_reg, col_reg}<16'b0110100100100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110100100100001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110100100100010) && ({row_reg, col_reg}<16'b0110100100100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110100100100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110100100100110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110100100100111) && ({row_reg, col_reg}<16'b0110100100101001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110100100101001) && ({row_reg, col_reg}<16'b0110100100101011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110100100101011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110100100101100) && ({row_reg, col_reg}<16'b0110100100101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110100100101110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110100100101111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110100100110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110100100110001) && ({row_reg, col_reg}<16'b0110100100110011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110100100110011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110100100110100) && ({row_reg, col_reg}<16'b0110100100111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110100100111010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110100100111011) && ({row_reg, col_reg}<16'b0110100101000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110100101000001) && ({row_reg, col_reg}<16'b0110100101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110100101000100) && ({row_reg, col_reg}<16'b0110100101001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110100101001001) && ({row_reg, col_reg}<16'b0110100101001100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110100101001100) && ({row_reg, col_reg}<16'b0110100101001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110100101001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110100101001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110100101010000) && ({row_reg, col_reg}<16'b0110100101011011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110100101011011) && ({row_reg, col_reg}<16'b0110100101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110100101011110) && ({row_reg, col_reg}<16'b0110100101100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110100101100001) && ({row_reg, col_reg}<16'b0110100101100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110100101100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100101100100) && ({row_reg, col_reg}<16'b0110100101101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110100101101000) && ({row_reg, col_reg}<16'b0110100101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100101101111) && ({row_reg, col_reg}<16'b0110100101110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100101110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100101110010) && ({row_reg, col_reg}<16'b0110100101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110100101110100) && ({row_reg, col_reg}<16'b0110100101111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100101111000) && ({row_reg, col_reg}<16'b0110100101111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100101111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110100101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100101111100) && ({row_reg, col_reg}<16'b0110100101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100101111110) && ({row_reg, col_reg}<16'b0110100110000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110100110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110100110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100110000011) && ({row_reg, col_reg}<16'b0110100110100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110100110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100110100101) && ({row_reg, col_reg}<16'b0110100110101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100110101000) && ({row_reg, col_reg}<16'b0110100110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100110101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110100110101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110100110101100) && ({row_reg, col_reg}<16'b0110100110101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110100110101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100110110000) && ({row_reg, col_reg}<16'b0110100110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110100110110110) && ({row_reg, col_reg}<16'b0110100110111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100110111010) && ({row_reg, col_reg}<16'b0110100110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100110111101) && ({row_reg, col_reg}<16'b0110100111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110100111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100111000001) && ({row_reg, col_reg}<16'b0110100111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110100111000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100111000100) && ({row_reg, col_reg}<16'b0110100111001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100111001111) && ({row_reg, col_reg}<16'b0110100111010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100111010001) && ({row_reg, col_reg}<16'b0110100111010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100111010011) && ({row_reg, col_reg}<16'b0110100111010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100111010110) && ({row_reg, col_reg}<16'b0110100111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100111011111) && ({row_reg, col_reg}<16'b0110100111100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110100111100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100111100010) && ({row_reg, col_reg}<16'b0110100111100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100111100111) && ({row_reg, col_reg}<16'b0110100111101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100111101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110100111101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100111101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110100111110000)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0110100111110001) && ({row_reg, col_reg}<16'b0110101000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110101000000000) && ({row_reg, col_reg}<16'b0110101000000100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110101000000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101000000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110101000000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110101000000111) && ({row_reg, col_reg}<16'b0110101000001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110101000001001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110101000001010) && ({row_reg, col_reg}<16'b0110101000001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101000001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110101000001101) && ({row_reg, col_reg}<16'b0110101000001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110101000001111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110101000010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101000010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110101000010010) && ({row_reg, col_reg}<16'b0110101000011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110101000011000) && ({row_reg, col_reg}<16'b0110101000011010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110101000011010) && ({row_reg, col_reg}<16'b0110101000011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110101000011100) && ({row_reg, col_reg}<16'b0110101000011110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110101000011110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110101000011111) && ({row_reg, col_reg}<16'b0110101000100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110101000100001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110101000100010) && ({row_reg, col_reg}<16'b0110101000100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110101000100101) && ({row_reg, col_reg}<16'b0110101000100111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110101000100111) && ({row_reg, col_reg}<16'b0110101000101010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110101000101010) && ({row_reg, col_reg}<16'b0110101000101100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110101000101100) && ({row_reg, col_reg}<16'b0110101000101110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110101000101110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110101000101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110101000110000) && ({row_reg, col_reg}<16'b0110101000110011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110101000110011) && ({row_reg, col_reg}<16'b0110101000110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110101000110111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110101000111000) && ({row_reg, col_reg}<16'b0110101001001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101001001001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110101001001010) && ({row_reg, col_reg}<16'b0110101001010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110101001010001) && ({row_reg, col_reg}<16'b0110101001010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110101001010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110101001010101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110101001010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110101001010111) && ({row_reg, col_reg}<16'b0110101001011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101001011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110101001011101) && ({row_reg, col_reg}<16'b0110101001011111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110101001011111) && ({row_reg, col_reg}<16'b0110101001100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110101001100001) && ({row_reg, col_reg}<16'b0110101001100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110101001100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110101001100101) && ({row_reg, col_reg}<16'b0110101001101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110101001101010) && ({row_reg, col_reg}<16'b0110101001110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110101001110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110101001110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101001110010) && ({row_reg, col_reg}<16'b0110101001110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110101001110100) && ({row_reg, col_reg}<16'b0110101001111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110101001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101001111001) && ({row_reg, col_reg}<16'b0110101001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110101001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101001111100) && ({row_reg, col_reg}<16'b0110101001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110101001111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110101010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110101010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101010000011) && ({row_reg, col_reg}<16'b0110101010100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110101010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101010100101) && ({row_reg, col_reg}<16'b0110101010101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110101010101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101010101001) && ({row_reg, col_reg}<16'b0110101010101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110101010101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110101010101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101010101101) && ({row_reg, col_reg}<16'b0110101010101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110101010101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101010110000) && ({row_reg, col_reg}<16'b0110101010110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110101010110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101010110110) && ({row_reg, col_reg}<16'b0110101010111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110101010111001) && ({row_reg, col_reg}<16'b0110101010111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101010111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110101010111100) && ({row_reg, col_reg}<16'b0110101010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101010111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110101010111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101011000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101011000001) && ({row_reg, col_reg}<16'b0110101011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110101011000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110101011000100) && ({row_reg, col_reg}<16'b0110101011001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101011001111) && ({row_reg, col_reg}<16'b0110101011010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110101011010001) && ({row_reg, col_reg}<16'b0110101011010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101011010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110101011010101) && ({row_reg, col_reg}<16'b0110101011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101011011111) && ({row_reg, col_reg}<16'b0110101011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110101011100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101011100010) && ({row_reg, col_reg}<16'b0110101011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110101011100111) && ({row_reg, col_reg}<16'b0110101011101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101011101001) && ({row_reg, col_reg}<16'b0110101011101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101011101100) && ({row_reg, col_reg}<16'b0110101011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101011101111) && ({row_reg, col_reg}<16'b0110101011110001)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0110101011110001) && ({row_reg, col_reg}<16'b0110101100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110101100000000) && ({row_reg, col_reg}<16'b0110101100000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110101100000100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110101100000101) && ({row_reg, col_reg}<16'b0110101100010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110101100010011) && ({row_reg, col_reg}<16'b0110101100010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110101100010101) && ({row_reg, col_reg}<16'b0110101100011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101100011011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110101100011100) && ({row_reg, col_reg}<16'b0110101100100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110101100100011) && ({row_reg, col_reg}<16'b0110101100101110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110101100101110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110101100101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110101100110000) && ({row_reg, col_reg}<16'b0110101100110100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110101100110100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110101100110101) && ({row_reg, col_reg}<16'b0110101101000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110101101000010) && ({row_reg, col_reg}<16'b0110101101000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110101101000100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110101101000101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110101101000110) && ({row_reg, col_reg}<16'b0110101101001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101101001001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110101101001010) && ({row_reg, col_reg}<16'b0110101101010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110101101010001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110101101010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101101010011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110101101010100) && ({row_reg, col_reg}<16'b0110101101010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110101101010110) && ({row_reg, col_reg}<16'b0110101101011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110101101011010) && ({row_reg, col_reg}<16'b0110101101011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110101101011100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0110101101011101) && ({row_reg, col_reg}<16'b0110101101011111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110101101011111) && ({row_reg, col_reg}<16'b0110101101101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110101101101011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0110101101101100) && ({row_reg, col_reg}<16'b0110101101101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110101101101110) && ({row_reg, col_reg}<16'b0110101101110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101101110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110101101110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101101110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110101101110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110101101110100) && ({row_reg, col_reg}<16'b0110101101111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110101101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101101111001) && ({row_reg, col_reg}<16'b0110101101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110101101111011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==16'b0110101101111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110101101111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101101111110) && ({row_reg, col_reg}<16'b0110101110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110101110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101110000011) && ({row_reg, col_reg}<16'b0110101110100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110101110100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101110100100) && ({row_reg, col_reg}<16'b0110101110100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110101110100111) && ({row_reg, col_reg}<16'b0110101110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101110101001) && ({row_reg, col_reg}<16'b0110101110101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110101110101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110101110101100) && ({row_reg, col_reg}<16'b0110101110101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110101110101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101110110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101110110001) && ({row_reg, col_reg}<16'b0110101110110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110101110110100) && ({row_reg, col_reg}<16'b0110101110110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101110110110) && ({row_reg, col_reg}<16'b0110101110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110101110111000) && ({row_reg, col_reg}<16'b0110101110111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101110111010) && ({row_reg, col_reg}<16'b0110101110111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110101110111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101111000000) && ({row_reg, col_reg}<16'b0110101111000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110101111000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101111000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110101111000100) && ({row_reg, col_reg}<16'b0110101111001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101111001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110101111001011) && ({row_reg, col_reg}<16'b0110101111001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101111001111) && ({row_reg, col_reg}<16'b0110101111010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110101111010001) && ({row_reg, col_reg}<16'b0110101111011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101111011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110101111011101) && ({row_reg, col_reg}<16'b0110101111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101111011111) && ({row_reg, col_reg}<16'b0110101111100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110101111100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101111100010) && ({row_reg, col_reg}<16'b0110101111100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110101111100111) && ({row_reg, col_reg}<16'b0110101111101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101111101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101111101010) && ({row_reg, col_reg}<16'b0110101111110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101111110000)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0110101111110001) && ({row_reg, col_reg}<16'b0110110000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110110000000000) && ({row_reg, col_reg}<16'b0110110000000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110110000000101) && ({row_reg, col_reg}<16'b0110110000011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110000011101)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0110110000011110) && ({row_reg, col_reg}<16'b0110110000100001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110110000100001) && ({row_reg, col_reg}<16'b0110110000100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110110000100110) && ({row_reg, col_reg}<16'b0110110000101010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110110000101010) && ({row_reg, col_reg}<16'b0110110000101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110110000101100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110110000101101) && ({row_reg, col_reg}<16'b0110110000110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110110000110010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110110000110011) && ({row_reg, col_reg}<16'b0110110000111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110110000111001) && ({row_reg, col_reg}<16'b0110110000111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110110000111011) && ({row_reg, col_reg}<16'b0110110001000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110001000001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110110001000010) && ({row_reg, col_reg}<16'b0110110001000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110110001000111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110110001001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110001001001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110110001001010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110110001001011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110110001001100) && ({row_reg, col_reg}<16'b0110110001010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110110001010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110110001010011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110110001010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110110001010101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110110001010110) && ({row_reg, col_reg}<16'b0110110001011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110001011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110110001011001) && ({row_reg, col_reg}<16'b0110110001011101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110110001011101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110110001011110) && ({row_reg, col_reg}<16'b0110110001101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110110001101000) && ({row_reg, col_reg}<16'b0110110001101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110001101011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0110110001101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110110001101101) && ({row_reg, col_reg}<16'b0110110001110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110001110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110110001110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110001110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110110001110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110110001110100) && ({row_reg, col_reg}<16'b0110110001111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110110001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110001111001) && ({row_reg, col_reg}<16'b0110110001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110110001111011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==16'b0110110001111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110001111101) && ({row_reg, col_reg}<16'b0110110001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110010000000) && ({row_reg, col_reg}<16'b0110110010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110010000011) && ({row_reg, col_reg}<16'b0110110010100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110010100100) && ({row_reg, col_reg}<16'b0110110010100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110010100111) && ({row_reg, col_reg}<16'b0110110010101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110010101001) && ({row_reg, col_reg}<16'b0110110010101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110010101011) && ({row_reg, col_reg}<16'b0110110010101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110110010101110) && ({row_reg, col_reg}<16'b0110110010110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110010110000) && ({row_reg, col_reg}<16'b0110110010110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110110010110100) && ({row_reg, col_reg}<16'b0110110010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110010110110) && ({row_reg, col_reg}<16'b0110110010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110010111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110110010111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110010111010) && ({row_reg, col_reg}<16'b0110110010111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110110010111111) && ({row_reg, col_reg}<16'b0110110011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110011000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110011000010) && ({row_reg, col_reg}<16'b0110110011000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110011000100) && ({row_reg, col_reg}<16'b0110110011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110011001011) && ({row_reg, col_reg}<16'b0110110011001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110011001111) && ({row_reg, col_reg}<16'b0110110011010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110011010001) && ({row_reg, col_reg}<16'b0110110011011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110011011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110110011011101) && ({row_reg, col_reg}<16'b0110110011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110011011111) && ({row_reg, col_reg}<16'b0110110011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110011100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110011100010) && ({row_reg, col_reg}<16'b0110110011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110011100111) && ({row_reg, col_reg}<16'b0110110011101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110011101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110011101010) && ({row_reg, col_reg}<16'b0110110011110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110011110000)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0110110011110001) && ({row_reg, col_reg}<16'b0110110100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110110100000000) && ({row_reg, col_reg}<16'b0110110100000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110110100000101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110110100000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110110100000111) && ({row_reg, col_reg}<16'b0110110100001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110110100001001) && ({row_reg, col_reg}<16'b0110110100001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110110100001011) && ({row_reg, col_reg}<16'b0110110100001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110110100001110) && ({row_reg, col_reg}<16'b0110110100011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110100011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110110100011011) && ({row_reg, col_reg}<16'b0110110100100100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110100100100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110110100100101) && ({row_reg, col_reg}<16'b0110110100101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110110100101101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110110100101110) && ({row_reg, col_reg}<16'b0110110100110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110110100110111) && ({row_reg, col_reg}<16'b0110110100111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110110100111101) && ({row_reg, col_reg}<16'b0110110101001000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110110101001000) && ({row_reg, col_reg}<16'b0110110101001010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110110101001010) && ({row_reg, col_reg}<16'b0110110101010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110110101010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110110101010011) && ({row_reg, col_reg}<16'b0110110101010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110110101010110) && ({row_reg, col_reg}<16'b0110110101011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110110101011001) && ({row_reg, col_reg}<16'b0110110101011011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110110101011011) && ({row_reg, col_reg}<16'b0110110101011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110110101011110) && ({row_reg, col_reg}<16'b0110110101100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110110101100111) && ({row_reg, col_reg}<16'b0110110101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110110101101010) && ({row_reg, col_reg}<16'b0110110101101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110110101101111) && ({row_reg, col_reg}<16'b0110110101110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110110101110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110101110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110110101110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110110101110100) && ({row_reg, col_reg}<16'b0110110101111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110101111000) && ({row_reg, col_reg}<16'b0110110101111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110101111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110110101111011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=16'b0110110101111100) && ({row_reg, col_reg}<16'b0110110110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110110000000) && ({row_reg, col_reg}<16'b0110110110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110110000011) && ({row_reg, col_reg}<16'b0110110110100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110110100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110110100100) && ({row_reg, col_reg}<16'b0110110110100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110110110100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110110100111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110110101000) && ({row_reg, col_reg}<16'b0110110110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110110101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110110101011) && ({row_reg, col_reg}<16'b0110110110101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110110101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110110110101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110110110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110110110001) && ({row_reg, col_reg}<16'b0110110110110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110110110110100) && ({row_reg, col_reg}<16'b0110110110110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110110110110) && ({row_reg, col_reg}<16'b0110110110111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110110111001) && ({row_reg, col_reg}<16'b0110110110111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110110111011) && ({row_reg, col_reg}<16'b0110110110111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110110110111110) && ({row_reg, col_reg}<16'b0110110111000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110111000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110111000011) && ({row_reg, col_reg}<16'b0110110111001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110111001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110111001011) && ({row_reg, col_reg}<16'b0110110111010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110111010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110111010001) && ({row_reg, col_reg}<16'b0110110111010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110111010110) && ({row_reg, col_reg}<16'b0110110111011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110111011010) && ({row_reg, col_reg}<16'b0110110111011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110111011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110110111011101) && ({row_reg, col_reg}<16'b0110110111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110111011111) && ({row_reg, col_reg}<16'b0110110111100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110111100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110111100010) && ({row_reg, col_reg}<16'b0110110111100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110111100111) && ({row_reg, col_reg}<16'b0110110111101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110111101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110110111101101) && ({row_reg, col_reg}<16'b0110110111110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110111110000)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0110110111110001) && ({row_reg, col_reg}<16'b0110111000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110111000000000) && ({row_reg, col_reg}<16'b0110111000000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111000000100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110111000000101) && ({row_reg, col_reg}<16'b0110111000000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110111000000111) && ({row_reg, col_reg}<16'b0110111000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111000001001) && ({row_reg, col_reg}<16'b0110111000001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110111000001011) && ({row_reg, col_reg}<16'b0110111000010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111000010000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110111000010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110111000010010) && ({row_reg, col_reg}<16'b0110111000010101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110111000010101) && ({row_reg, col_reg}<16'b0110111000010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111000010111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110111000011000) && ({row_reg, col_reg}<16'b0110111000011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110111000011111) && ({row_reg, col_reg}<16'b0110111000100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111000100010) && ({row_reg, col_reg}<16'b0110111000100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110111000100111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0110111000101000) && ({row_reg, col_reg}<16'b0110111000101010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110111000101010) && ({row_reg, col_reg}<16'b0110111000111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110111000111000) && ({row_reg, col_reg}<16'b0110111000111100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110111000111100) && ({row_reg, col_reg}<16'b0110111001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111001001001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110111001001010) && ({row_reg, col_reg}<16'b0110111001010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111001010000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110111001010001) && ({row_reg, col_reg}<16'b0110111001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110111001010100) && ({row_reg, col_reg}<16'b0110111001011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111001011011) && ({row_reg, col_reg}<16'b0110111001100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110111001100111) && ({row_reg, col_reg}<16'b0110111001110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110111001110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110111001110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111001110010) && ({row_reg, col_reg}<16'b0110111001110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110111001110110) && ({row_reg, col_reg}<16'b0110111001111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111001111000) && ({row_reg, col_reg}<16'b0110111001111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111001111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111001111011) && ({row_reg, col_reg}<16'b0110111001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110111001111101) && ({row_reg, col_reg}<16'b0110111001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110111001111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110111010000000) && ({row_reg, col_reg}<16'b0110111010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111010000011) && ({row_reg, col_reg}<16'b0110111010100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110111010100100) && ({row_reg, col_reg}<16'b0110111010100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111010100110) && ({row_reg, col_reg}<16'b0110111010101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111010101000) && ({row_reg, col_reg}<16'b0110111010101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111010101011) && ({row_reg, col_reg}<16'b0110111010101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110111010101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111010101111) && ({row_reg, col_reg}<16'b0110111010110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111010110001) && ({row_reg, col_reg}<16'b0110111010110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110111010110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110111010110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111010110110) && ({row_reg, col_reg}<16'b0110111010111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111010111001) && ({row_reg, col_reg}<16'b0110111011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111011000001) && ({row_reg, col_reg}<16'b0110111011000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111011000011) && ({row_reg, col_reg}<16'b0110111011001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111011001100) && ({row_reg, col_reg}<16'b0110111011010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111011010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111011010001) && ({row_reg, col_reg}<16'b0110111011010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111011010101) && ({row_reg, col_reg}<16'b0110111011011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111011011010) && ({row_reg, col_reg}<16'b0110111011011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111011011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110111011011101) && ({row_reg, col_reg}<16'b0110111011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111011011111) && ({row_reg, col_reg}<16'b0110111011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110111011100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111011100010) && ({row_reg, col_reg}<16'b0110111011100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111011100100) && ({row_reg, col_reg}<16'b0110111011110001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0110111011110001) && ({row_reg, col_reg}<16'b0110111100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110111100000000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110111100000001) && ({row_reg, col_reg}<16'b0110111100000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111100000011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110111100000100) && ({row_reg, col_reg}<16'b0110111100000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110111100000110) && ({row_reg, col_reg}<16'b0110111100001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111100001001) && ({row_reg, col_reg}<16'b0110111100001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110111100001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111100001100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110111100001101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110111100001110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110111100001111) && ({row_reg, col_reg}<16'b0110111100011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111100011000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110111100011001) && ({row_reg, col_reg}<16'b0110111100011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110111100011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110111100011101) && ({row_reg, col_reg}<16'b0110111100100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110111100100000) && ({row_reg, col_reg}<16'b0110111100100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111100100010) && ({row_reg, col_reg}<16'b0110111100110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110111100110111) && ({row_reg, col_reg}<16'b0110111101001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111101001111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110111101010000) && ({row_reg, col_reg}<16'b0110111101010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110111101010010) && ({row_reg, col_reg}<16'b0110111101011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111101011000) && ({row_reg, col_reg}<16'b0110111101100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110111101100111) && ({row_reg, col_reg}<16'b0110111101101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111101101001) && ({row_reg, col_reg}<16'b0110111101101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0110111101101011) && ({row_reg, col_reg}<16'b0110111101101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111101101101) && ({row_reg, col_reg}<16'b0110111101110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110111101110000) && ({row_reg, col_reg}<16'b0110111101110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111101110010) && ({row_reg, col_reg}<16'b0110111101111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110111101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111101111001) && ({row_reg, col_reg}<16'b0110111101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110111101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111101111100) && ({row_reg, col_reg}<16'b0110111110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111110000000) && ({row_reg, col_reg}<16'b0110111110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111110000010) && ({row_reg, col_reg}<16'b0110111110100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110111110100100) && ({row_reg, col_reg}<16'b0110111110100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111110100110) && ({row_reg, col_reg}<16'b0110111110101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111110101000) && ({row_reg, col_reg}<16'b0110111110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111110101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111110101100) && ({row_reg, col_reg}<16'b0110111110101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110111110101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111110101111) && ({row_reg, col_reg}<16'b0110111110110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111110110001) && ({row_reg, col_reg}<16'b0110111110110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110111110110100) && ({row_reg, col_reg}<16'b0110111110110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111110110110) && ({row_reg, col_reg}<16'b0110111110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110111110111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111110111001) && ({row_reg, col_reg}<16'b0110111111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111111000000) && ({row_reg, col_reg}<16'b0110111111000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111111000011) && ({row_reg, col_reg}<16'b0110111111000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111111000110) && ({row_reg, col_reg}<16'b0110111111001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111111001000) && ({row_reg, col_reg}<16'b0110111111001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111111001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111111001101) && ({row_reg, col_reg}<16'b0110111111010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111111010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111111010001) && ({row_reg, col_reg}<16'b0110111111010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111111010110) && ({row_reg, col_reg}<16'b0110111111011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111111011010) && ({row_reg, col_reg}<16'b0110111111011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111111011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110111111011101) && ({row_reg, col_reg}<16'b0110111111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111111011111) && ({row_reg, col_reg}<16'b0110111111100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110111111100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111111100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111111100011) && ({row_reg, col_reg}<16'b0110111111101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111111101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111111101110) && ({row_reg, col_reg}<16'b0110111111110001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0110111111110001) && ({row_reg, col_reg}<16'b0111000000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000000000000) && ({row_reg, col_reg}<16'b0111000000000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111000000000010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111000000000011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111000000000100) && ({row_reg, col_reg}<16'b0111000000000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111000000000110) && ({row_reg, col_reg}<16'b0111000000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000000001001) && ({row_reg, col_reg}<16'b0111000000001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111000000001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111000000001100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111000000001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111000000001110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111000000001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111000000010000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111000000010001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111000000010010) && ({row_reg, col_reg}<16'b0111000000011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111000000011000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111000000011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111000000011010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111000000011011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111000000011100) && ({row_reg, col_reg}<16'b0111000000011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111000000011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111000000011111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111000000100000) && ({row_reg, col_reg}<16'b0111000000110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111000000110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111000000110011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111000000110100) && ({row_reg, col_reg}<16'b0111000000110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111000000110110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111000000110111) && ({row_reg, col_reg}<16'b0111000000111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111000000111100) && ({row_reg, col_reg}<16'b0111000001000000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111000001000000) && ({row_reg, col_reg}<16'b0111000001001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111000001001100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111000001001101) && ({row_reg, col_reg}<16'b0111000001010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111000001010001) && ({row_reg, col_reg}<16'b0111000001010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111000001010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111000001010100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0111000001010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000001010110) && ({row_reg, col_reg}<16'b0111000001101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111000001101000) && ({row_reg, col_reg}<16'b0111000001101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000001101100) && ({row_reg, col_reg}<16'b0111000001101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111000001101111) && ({row_reg, col_reg}<16'b0111000001111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000001111001) && ({row_reg, col_reg}<16'b0111000001111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000001111111) && ({row_reg, col_reg}<16'b0111000010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111000010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000010000010) && ({row_reg, col_reg}<16'b0111000010100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000010100011) && ({row_reg, col_reg}<16'b0111000010100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111000010100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000010100110) && ({row_reg, col_reg}<16'b0111000010101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000010101001) && ({row_reg, col_reg}<16'b0111000010101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000010101100) && ({row_reg, col_reg}<16'b0111000010101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111000010101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000010101111) && ({row_reg, col_reg}<16'b0111000010110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000010110001) && ({row_reg, col_reg}<16'b0111000010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111000010110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000010110100) && ({row_reg, col_reg}<16'b0111000010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111000010110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000010110111) && ({row_reg, col_reg}<16'b0111000010111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000010111001) && ({row_reg, col_reg}<16'b0111000011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000011000000) && ({row_reg, col_reg}<16'b0111000011000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000011000011) && ({row_reg, col_reg}<16'b0111000011000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000011000110) && ({row_reg, col_reg}<16'b0111000011001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000011001000) && ({row_reg, col_reg}<16'b0111000011001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000011001111) && ({row_reg, col_reg}<16'b0111000011010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000011010001) && ({row_reg, col_reg}<16'b0111000011010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000011010111) && ({row_reg, col_reg}<16'b0111000011011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000011011010) && ({row_reg, col_reg}<16'b0111000011011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111000011011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111000011011101) && ({row_reg, col_reg}<16'b0111000011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000011011111) && ({row_reg, col_reg}<16'b0111000011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000011100001) && ({row_reg, col_reg}<16'b0111000011101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111000011101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000011101110) && ({row_reg, col_reg}<16'b0111000011110001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0111000011110001) && ({row_reg, col_reg}<16'b0111000100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111000100000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000100000001) && ({row_reg, col_reg}<16'b0111000100000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111000100000101) && ({row_reg, col_reg}<16'b0111000100001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000100001001) && ({row_reg, col_reg}<16'b0111000100001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111000100001011) && ({row_reg, col_reg}<16'b0111000100001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111000100001101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111000100001110) && ({row_reg, col_reg}<16'b0111000100010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111000100010000) && ({row_reg, col_reg}<16'b0111000100010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111000100010010) && ({row_reg, col_reg}<16'b0111000100011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111000100011000) && ({row_reg, col_reg}<16'b0111000100011011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111000100011011) && ({row_reg, col_reg}<16'b0111000100100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111000100100010) && ({row_reg, col_reg}<16'b0111000100100100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111000100100100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111000100100101) && ({row_reg, col_reg}<16'b0111000100101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111000100101100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111000100101101) && ({row_reg, col_reg}<16'b0111000100110000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111000100110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111000100110001) && ({row_reg, col_reg}<16'b0111000100110100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111000100110100) && ({row_reg, col_reg}<16'b0111000100110111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111000100110111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111000100111000) && ({row_reg, col_reg}<16'b0111000100111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111000100111011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111000100111100) && ({row_reg, col_reg}<16'b0111000100111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111000100111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111000101000000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111000101000001) && ({row_reg, col_reg}<16'b0111000101001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111000101001011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111000101001100) && ({row_reg, col_reg}<16'b0111000101001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111000101001110) && ({row_reg, col_reg}<16'b0111000101010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000101010101) && ({row_reg, col_reg}<16'b0111000101100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111000101100001) && ({row_reg, col_reg}<16'b0111000101100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000101100100) && ({row_reg, col_reg}<16'b0111000101101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111000101101001) && ({row_reg, col_reg}<16'b0111000101101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111000101101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111000101101100) && ({row_reg, col_reg}<16'b0111000101101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000101101111) && ({row_reg, col_reg}<16'b0111000101110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111000101110001) && ({row_reg, col_reg}<16'b0111000101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000101111000) && ({row_reg, col_reg}<16'b0111000110000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111000110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000110000010) && ({row_reg, col_reg}<16'b0111000110100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000110100010) && ({row_reg, col_reg}<16'b0111000110100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111000110100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000110100110) && ({row_reg, col_reg}<16'b0111000110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000110101001) && ({row_reg, col_reg}<16'b0111000110101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111000110101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111000110101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000110101110) && ({row_reg, col_reg}<16'b0111000110110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000110110000) && ({row_reg, col_reg}<16'b0111000110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000110110011) && ({row_reg, col_reg}<16'b0111000110110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111000110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000110110111) && ({row_reg, col_reg}<16'b0111000110111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000110111010) && ({row_reg, col_reg}<16'b0111000111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000111000001) && ({row_reg, col_reg}<16'b0111000111000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000111000100) && ({row_reg, col_reg}<16'b0111000111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111000111000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000111001000) && ({row_reg, col_reg}<16'b0111000111001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000111001111) && ({row_reg, col_reg}<16'b0111000111010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000111010001) && ({row_reg, col_reg}<16'b0111000111010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000111010111) && ({row_reg, col_reg}<16'b0111000111011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000111011010) && ({row_reg, col_reg}<16'b0111000111011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111000111011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111000111011101) && ({row_reg, col_reg}<16'b0111000111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000111011111) && ({row_reg, col_reg}<16'b0111000111100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111000111100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000111100010) && ({row_reg, col_reg}<16'b0111000111110001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0111000111110001) && ({row_reg, col_reg}<16'b0111001000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001000000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001000000001) && ({row_reg, col_reg}<16'b0111001000000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111001000000011) && ({row_reg, col_reg}<16'b0111001000000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001000000111) && ({row_reg, col_reg}<16'b0111001000001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001000001010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0111001000001011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111001000001100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0111001000001101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111001000001110) && ({row_reg, col_reg}<16'b0111001000010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001000010000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111001000010001) && ({row_reg, col_reg}<16'b0111001000011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111001000011101) && ({row_reg, col_reg}<16'b0111001000011111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111001000011111) && ({row_reg, col_reg}<16'b0111001000100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111001000100110) && ({row_reg, col_reg}<16'b0111001000101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001000101010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111001000101011) && ({row_reg, col_reg}<16'b0111001000110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111001000110101) && ({row_reg, col_reg}<16'b0111001000110111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111001000110111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111001000111000) && ({row_reg, col_reg}<16'b0111001000111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111001000111100) && ({row_reg, col_reg}<16'b0111001000111110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111001000111110) && ({row_reg, col_reg}<16'b0111001001000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001001000100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111001001000101) && ({row_reg, col_reg}<16'b0111001001000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111001001000111) && ({row_reg, col_reg}<16'b0111001001001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001001001001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111001001001010) && ({row_reg, col_reg}<16'b0111001001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111001001001100) && ({row_reg, col_reg}<16'b0111001001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111001001001110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0111001001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001001010000) && ({row_reg, col_reg}<16'b0111001001011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001001011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111001001011110) && ({row_reg, col_reg}<16'b0111001001100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111001001100001) && ({row_reg, col_reg}<16'b0111001001100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001001100100) && ({row_reg, col_reg}<16'b0111001001101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001001101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001001101010) && ({row_reg, col_reg}<16'b0111001001101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111001001101100) && ({row_reg, col_reg}<16'b0111001001101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001001101110) && ({row_reg, col_reg}<16'b0111001001110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001001110000) && ({row_reg, col_reg}<16'b0111001001110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001001110010) && ({row_reg, col_reg}<16'b0111001001110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111001001110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001001110110) && ({row_reg, col_reg}<16'b0111001010000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111001010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001010000010) && ({row_reg, col_reg}<16'b0111001010100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001010100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001010100010) && ({row_reg, col_reg}<16'b0111001010100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001010100101) && ({row_reg, col_reg}<16'b0111001010101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001010101000) && ({row_reg, col_reg}<16'b0111001010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001010101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111001010101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001010101100) && ({row_reg, col_reg}<16'b0111001010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001010110000) && ({row_reg, col_reg}<16'b0111001010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001010110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001010110100) && ({row_reg, col_reg}<16'b0111001010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001010110110) && ({row_reg, col_reg}<16'b0111001010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111001010111000) && ({row_reg, col_reg}<16'b0111001010111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001010111010) && ({row_reg, col_reg}<16'b0111001010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001010111100) && ({row_reg, col_reg}<16'b0111001011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001011000001) && ({row_reg, col_reg}<16'b0111001011000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001011000100) && ({row_reg, col_reg}<16'b0111001011010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001011010110) && ({row_reg, col_reg}<16'b0111001011011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001011011010) && ({row_reg, col_reg}<16'b0111001011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001011011111) && ({row_reg, col_reg}<16'b0111001011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001011100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111001011100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001011100011) && ({row_reg, col_reg}<16'b0111001011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001011100111) && ({row_reg, col_reg}<16'b0111001011101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001011101110) && ({row_reg, col_reg}<16'b0111001011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111001011110000)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0111001011110001) && ({row_reg, col_reg}<16'b0111001100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001100000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001100000001) && ({row_reg, col_reg}<16'b0111001100000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001100000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111001100000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111001100000101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0111001100000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001100000111) && ({row_reg, col_reg}<16'b0111001100001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001100001010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111001100001011)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0111001100001100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111001100001101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111001100001110) && ({row_reg, col_reg}<16'b0111001100011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111001100011101) && ({row_reg, col_reg}<16'b0111001100011111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111001100011111) && ({row_reg, col_reg}<16'b0111001100100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001100100110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111001100100111) && ({row_reg, col_reg}<16'b0111001100101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111001100101001) && ({row_reg, col_reg}<16'b0111001100101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111001100101101) && ({row_reg, col_reg}<16'b0111001100101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111001100101111) && ({row_reg, col_reg}<16'b0111001100110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001100110101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111001100110110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111001100110111) && ({row_reg, col_reg}<16'b0111001101001000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111001101001000) && ({row_reg, col_reg}<16'b0111001101001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001101001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001101001011) && ({row_reg, col_reg}<16'b0111001101001101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0111001101001101) && ({row_reg, col_reg}<16'b0111001101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001101001111) && ({row_reg, col_reg}<16'b0111001101011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111001101011001) && ({row_reg, col_reg}<16'b0111001101011011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111001101011011) && ({row_reg, col_reg}<16'b0111001101100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111001101100111) && ({row_reg, col_reg}<16'b0111001101101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111001101101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111001101101010) && ({row_reg, col_reg}<16'b0111001101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001101101110) && ({row_reg, col_reg}<16'b0111001110000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111001110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001110000011) && ({row_reg, col_reg}<16'b0111001110100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001110100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001110100010) && ({row_reg, col_reg}<16'b0111001110100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111001110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001110100101) && ({row_reg, col_reg}<16'b0111001110100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001110100111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001110101000) && ({row_reg, col_reg}<16'b0111001110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001110101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001110101011) && ({row_reg, col_reg}<16'b0111001110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001110110000) && ({row_reg, col_reg}<16'b0111001110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001110110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111001110110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001110110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001110110110) && ({row_reg, col_reg}<16'b0111001110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111001110111000) && ({row_reg, col_reg}<16'b0111001110111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001110111100) && ({row_reg, col_reg}<16'b0111001111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001111000001) && ({row_reg, col_reg}<16'b0111001111000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001111000011) && ({row_reg, col_reg}<16'b0111001111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001111000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001111000110) && ({row_reg, col_reg}<16'b0111001111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001111001000) && ({row_reg, col_reg}<16'b0111001111001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001111001010) && ({row_reg, col_reg}<16'b0111001111010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001111010101) && ({row_reg, col_reg}<16'b0111001111011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001111011010) && ({row_reg, col_reg}<16'b0111001111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001111011111) && ({row_reg, col_reg}<16'b0111001111100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001111100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001111100010) && ({row_reg, col_reg}<16'b0111001111100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001111100111) && ({row_reg, col_reg}<16'b0111001111101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001111101110) && ({row_reg, col_reg}<16'b0111001111110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111001111110000)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b0111001111110001) && ({row_reg, col_reg}<16'b0111010000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111010000000000) && ({row_reg, col_reg}<16'b0111010000000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111010000000100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0111010000000101) && ({row_reg, col_reg}<16'b0111010000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111010000001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111010000001010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111010000001011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111010000001100) && ({row_reg, col_reg}<16'b0111010000001110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111010000001110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111010000001111) && ({row_reg, col_reg}<16'b0111010000100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111010000100110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111010000100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111010000101000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111010000101001) && ({row_reg, col_reg}<16'b0111010000101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111010000101100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111010000101101) && ({row_reg, col_reg}<16'b0111010000101111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111010000101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111010000110000) && ({row_reg, col_reg}<16'b0111010001000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111010001000100) && ({row_reg, col_reg}<16'b0111010001000110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111010001000110) && ({row_reg, col_reg}<16'b0111010001001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111010001001001) && ({row_reg, col_reg}<16'b0111010001001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111010001001110) && ({row_reg, col_reg}<16'b0111010001010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111010001010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111010001010100) && ({row_reg, col_reg}<16'b0111010001011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111010001011001) && ({row_reg, col_reg}<16'b0111010001011011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111010001011011) && ({row_reg, col_reg}<16'b0111010001100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111010001100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111010001100111) && ({row_reg, col_reg}<16'b0111010001101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111010001101010) && ({row_reg, col_reg}<16'b0111010001101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010001101101) && ({row_reg, col_reg}<16'b0111010001110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111010001110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111010001110001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111010001110010) && ({row_reg, col_reg}<16'b0111010001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111010001111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111010001111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111010001111101) && ({row_reg, col_reg}<16'b0111010001111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111010001111111) && ({row_reg, col_reg}<16'b0111010010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010010000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010010000011) && ({row_reg, col_reg}<16'b0111010010011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111010010011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010010011110) && ({row_reg, col_reg}<16'b0111010010100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111010010100010) && ({row_reg, col_reg}<16'b0111010010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010010100100) && ({row_reg, col_reg}<16'b0111010010101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111010010101000) && ({row_reg, col_reg}<16'b0111010010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010010101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010010101011) && ({row_reg, col_reg}<16'b0111010010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111010010110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010010110001) && ({row_reg, col_reg}<16'b0111010010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111010010110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111010010110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010010110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010010110110) && ({row_reg, col_reg}<16'b0111010010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111010010111000) && ({row_reg, col_reg}<16'b0111010010111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111010010111011) && ({row_reg, col_reg}<16'b0111010011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010011000000) && ({row_reg, col_reg}<16'b0111010011000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111010011000011) && ({row_reg, col_reg}<16'b0111010011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010011001001) && ({row_reg, col_reg}<16'b0111010011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111010011001011) && ({row_reg, col_reg}<16'b0111010011010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010011010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111010011010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010011010101) && ({row_reg, col_reg}<16'b0111010011010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111010011010111) && ({row_reg, col_reg}<16'b0111010011011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010011011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111010011011010) && ({row_reg, col_reg}<16'b0111010011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010011011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111010011100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010011100001) && ({row_reg, col_reg}<16'b0111010011100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010011100011) && ({row_reg, col_reg}<16'b0111010011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111010011100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010011101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010011101001) && ({row_reg, col_reg}<16'b0111010011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010011101111) && ({row_reg, col_reg}<16'b0111010011110001)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0111010011110001) && ({row_reg, col_reg}<16'b0111010100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111010100000000) && ({row_reg, col_reg}<16'b0111010100000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111010100000101) && ({row_reg, col_reg}<16'b0111010100001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111010100001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111010100001010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111010100001011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111010100001100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0111010100001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0111010100001110) && ({row_reg, col_reg}<16'b0111010100010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111010100010000) && ({row_reg, col_reg}<16'b0111010100010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111010100010010) && ({row_reg, col_reg}<16'b0111010100100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111010100100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111010100101000) && ({row_reg, col_reg}<16'b0111010100101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111010100101101) && ({row_reg, col_reg}<16'b0111010100110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111010100110000) && ({row_reg, col_reg}<16'b0111010101000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111010101000000) && ({row_reg, col_reg}<16'b0111010101000010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111010101000010) && ({row_reg, col_reg}<16'b0111010101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111010101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111010101000111) && ({row_reg, col_reg}<16'b0111010101001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111010101001001) && ({row_reg, col_reg}<16'b0111010101001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111010101001100) && ({row_reg, col_reg}<16'b0111010101100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111010101100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111010101100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111010101100111) && ({row_reg, col_reg}<16'b0111010101101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010101101100) && ({row_reg, col_reg}<16'b0111010101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111010101101111) && ({row_reg, col_reg}<16'b0111010101110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0111010101110010) && ({row_reg, col_reg}<16'b0111010101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111010101111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111010101111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111010101111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111010101111110) && ({row_reg, col_reg}<16'b0111010110000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010110000011) && ({row_reg, col_reg}<16'b0111010110000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010110000110) && ({row_reg, col_reg}<16'b0111010110001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010110001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111010110001100) && ({row_reg, col_reg}<16'b0111010110001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010110001110) && ({row_reg, col_reg}<16'b0111010110010111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010110010111) && ({row_reg, col_reg}<16'b0111010110011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010110011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010110011110) && ({row_reg, col_reg}<16'b0111010110101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111010110101000) && ({row_reg, col_reg}<16'b0111010110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010110101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010110101011) && ({row_reg, col_reg}<16'b0111010110101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111010110101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010110110000) && ({row_reg, col_reg}<16'b0111010110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111010110110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111010110110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010110110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010110110110) && ({row_reg, col_reg}<16'b0111010110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111010110111000) && ({row_reg, col_reg}<16'b0111010110111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111010110111010) && ({row_reg, col_reg}<16'b0111010110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010110111101) && ({row_reg, col_reg}<16'b0111010110111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010110111111) && ({row_reg, col_reg}<16'b0111010111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010111001000) && ({row_reg, col_reg}<16'b0111010111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111010111001011) && ({row_reg, col_reg}<16'b0111010111010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010111010100) && ({row_reg, col_reg}<16'b0111010111010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111010111010110) && ({row_reg, col_reg}<16'b0111010111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010111011111) && ({row_reg, col_reg}<16'b0111010111100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010111100001) && ({row_reg, col_reg}<16'b0111010111100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010111100011) && ({row_reg, col_reg}<16'b0111010111101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111010111101000) && ({row_reg, col_reg}<16'b0111010111101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010111101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111010111101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010111101111) && ({row_reg, col_reg}<16'b0111010111110001)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0111010111110001) && ({row_reg, col_reg}<16'b0111011000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111011000000000) && ({row_reg, col_reg}<16'b0111011000000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111011000000111) && ({row_reg, col_reg}<16'b0111011000001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111011000001001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111011000001010)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0111011000001011) && ({row_reg, col_reg}<16'b0111011000001101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0111011000001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111011000001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111011000001111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0111011000010000) && ({row_reg, col_reg}<16'b0111011000010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111011000010010) && ({row_reg, col_reg}<16'b0111011000010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111011000010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111011000010101) && ({row_reg, col_reg}<16'b0111011000111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111011000111111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111011001000000) && ({row_reg, col_reg}<16'b0111011001000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111011001000011) && ({row_reg, col_reg}<16'b0111011001000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111011001000101) && ({row_reg, col_reg}<16'b0111011001001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111011001001000) && ({row_reg, col_reg}<16'b0111011001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111011001001011) && ({row_reg, col_reg}<16'b0111011001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111011001011111) && ({row_reg, col_reg}<16'b0111011001100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111011001100001) && ({row_reg, col_reg}<16'b0111011001100100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111011001100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111011001100101) && ({row_reg, col_reg}<16'b0111011001100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111011001100111) && ({row_reg, col_reg}<16'b0111011001101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011001101001) && ({row_reg, col_reg}<16'b0111011001101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111011001101100) && ({row_reg, col_reg}<16'b0111011001101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011001101110) && ({row_reg, col_reg}<16'b0111011001110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111011001110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111011001110101) && ({row_reg, col_reg}<16'b0111011001110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011001110111) && ({row_reg, col_reg}<16'b0111011001111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111011001111001) && ({row_reg, col_reg}<16'b0111011001111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011001111101) && ({row_reg, col_reg}<16'b0111011010010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011010010111) && ({row_reg, col_reg}<16'b0111011010011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011010011001) && ({row_reg, col_reg}<16'b0111011010011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011010011100) && ({row_reg, col_reg}<16'b0111011010011110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011010011110) && ({row_reg, col_reg}<16'b0111011010100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111011010100111) && ({row_reg, col_reg}<16'b0111011010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011010101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111011010101011) && ({row_reg, col_reg}<16'b0111011010101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011010101110) && ({row_reg, col_reg}<16'b0111011010110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011010110000) && ({row_reg, col_reg}<16'b0111011010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111011010110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111011010110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011010110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011010110110) && ({row_reg, col_reg}<16'b0111011010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111011010111000) && ({row_reg, col_reg}<16'b0111011010111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011010111010) && ({row_reg, col_reg}<16'b0111011011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011011001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011011001001) && ({row_reg, col_reg}<16'b0111011011010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011011010100) && ({row_reg, col_reg}<16'b0111011011010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011011010111) && ({row_reg, col_reg}<16'b0111011011100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011011100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011011100001) && ({row_reg, col_reg}<16'b0111011011100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011011100011) && ({row_reg, col_reg}<16'b0111011011100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011011100110) && ({row_reg, col_reg}<16'b0111011011101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111011011101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111011011101011) && ({row_reg, col_reg}<16'b0111011011101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011011101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011011101110) && ({row_reg, col_reg}<16'b0111011011110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011011110000)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b0111011011110001) && ({row_reg, col_reg}<16'b0111011100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111011100000000) && ({row_reg, col_reg}<16'b0111011100000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111011100000101)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0111011100000110) && ({row_reg, col_reg}<16'b0111011100001010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111011100001010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111011100001011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0111011100001100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111011100001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111011100001110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0111011100001111) && ({row_reg, col_reg}<16'b0111011100010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111011100010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111011100010010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0111011100010011) && ({row_reg, col_reg}<16'b0111011100011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111011100011000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111011100011001) && ({row_reg, col_reg}<16'b0111011100110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111011100110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111011100110110) && ({row_reg, col_reg}<16'b0111011100111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111011100111110) && ({row_reg, col_reg}<16'b0111011101000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111011101000010) && ({row_reg, col_reg}<16'b0111011101000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111011101000100) && ({row_reg, col_reg}<16'b0111011101001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111011101001000) && ({row_reg, col_reg}<16'b0111011101100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111011101100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111011101100100) && ({row_reg, col_reg}<16'b0111011101101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111011101101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011101101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011101101010) && ({row_reg, col_reg}<16'b0111011101101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111011101101100) && ({row_reg, col_reg}<16'b0111011101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011101101110)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b0111011101101111) && ({row_reg, col_reg}<16'b0111011101110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111011101110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011101110101)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==16'b0111011101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011101110111) && ({row_reg, col_reg}<16'b0111011101111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111011101111001) && ({row_reg, col_reg}<16'b0111011101111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011101111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011101111110) && ({row_reg, col_reg}<16'b0111011110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011110000000) && ({row_reg, col_reg}<16'b0111011110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011110000010) && ({row_reg, col_reg}<16'b0111011110000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011110000100) && ({row_reg, col_reg}<16'b0111011110010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011110010011) && ({row_reg, col_reg}<16'b0111011110010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011110010101) && ({row_reg, col_reg}<16'b0111011110010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011110011000) && ({row_reg, col_reg}<16'b0111011110011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011110011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011110011110) && ({row_reg, col_reg}<16'b0111011110100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111011110100111) && ({row_reg, col_reg}<16'b0111011110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011110101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011110101011) && ({row_reg, col_reg}<16'b0111011110101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011110101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011110101111) && ({row_reg, col_reg}<16'b0111011110110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011110110001) && ({row_reg, col_reg}<16'b0111011110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111011110110011) && ({row_reg, col_reg}<16'b0111011110110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011110110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011110110110) && ({row_reg, col_reg}<16'b0111011110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111011110111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011110111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011110111010) && ({row_reg, col_reg}<16'b0111011111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011111001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011111001001) && ({row_reg, col_reg}<16'b0111011111001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011111001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011111001101) && ({row_reg, col_reg}<16'b0111011111010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011111010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011111010101) && ({row_reg, col_reg}<16'b0111011111100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011111100011) && ({row_reg, col_reg}<16'b0111011111100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011111100101) && ({row_reg, col_reg}<16'b0111011111100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111011111100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111011111101000) && ({row_reg, col_reg}<16'b0111011111101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111011111101010) && ({row_reg, col_reg}<16'b0111011111101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111011111101100) && ({row_reg, col_reg}<16'b0111011111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011111101111) && ({row_reg, col_reg}<16'b0111011111110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011111110001)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0111011111110010) && ({row_reg, col_reg}<16'b0111100000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111100000000000) && ({row_reg, col_reg}<16'b0111100000000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111100000000101) && ({row_reg, col_reg}<16'b0111100000001011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0111100000001011) && ({row_reg, col_reg}<16'b0111100000001101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111100000001101) && ({row_reg, col_reg}<16'b0111100000001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111100000001111) && ({row_reg, col_reg}<16'b0111100000011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111100000011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111100000011001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111100000011010) && ({row_reg, col_reg}<16'b0111100000111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111100000111100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111100000111101) && ({row_reg, col_reg}<16'b0111100000111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111100000111111) && ({row_reg, col_reg}<16'b0111100001000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111100001000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111100001000101) && ({row_reg, col_reg}<16'b0111100001000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111100001000111) && ({row_reg, col_reg}<16'b0111100001001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111100001001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111100001001110) && ({row_reg, col_reg}<16'b0111100001100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111100001100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111100001100010) && ({row_reg, col_reg}<16'b0111100001100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111100001100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111100001101000) && ({row_reg, col_reg}<16'b0111100001101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100001101010) && ({row_reg, col_reg}<16'b0111100001101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111100001101100) && ({row_reg, col_reg}<16'b0111100001110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100001110000) && ({row_reg, col_reg}<16'b0111100001110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0111100001110011) && ({row_reg, col_reg}<16'b0111100001110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111100001110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111100001110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0111100001110111) && ({row_reg, col_reg}<16'b0111100001111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111100001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100001111101) && ({row_reg, col_reg}<16'b0111100010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111100010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100010000001) && ({row_reg, col_reg}<16'b0111100010000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100010000100) && ({row_reg, col_reg}<16'b0111100010010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100010010010) && ({row_reg, col_reg}<16'b0111100010010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111100010010101) && ({row_reg, col_reg}<16'b0111100010011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100010011110) && ({row_reg, col_reg}<16'b0111100010100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111100010100001) && ({row_reg, col_reg}<16'b0111100010100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111100010100011) && ({row_reg, col_reg}<16'b0111100010100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111100010100111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111100010101000) && ({row_reg, col_reg}<16'b0111100010110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111100010110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111100010110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111100010110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111100010111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111100010111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100010111010) && ({row_reg, col_reg}<16'b0111100010111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100010111111) && ({row_reg, col_reg}<16'b0111100011000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100011000010) && ({row_reg, col_reg}<16'b0111100011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100011001001) && ({row_reg, col_reg}<16'b0111100011001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100011001101) && ({row_reg, col_reg}<16'b0111100011010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111100011010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100011010001) && ({row_reg, col_reg}<16'b0111100011100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100011100101) && ({row_reg, col_reg}<16'b0111100011100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111100011100111) && ({row_reg, col_reg}<16'b0111100011101001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111100011101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100011101010) && ({row_reg, col_reg}<16'b0111100011101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111100011101110) && ({row_reg, col_reg}<16'b0111100011110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111100011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111100011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111100011110010)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0111100011110011) && ({row_reg, col_reg}<16'b0111100100000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111100100000000) && ({row_reg, col_reg}<16'b0111100100000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111100100000101) && ({row_reg, col_reg}<16'b0111100100001001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0111100100001001) && ({row_reg, col_reg}<16'b0111100100001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111100100001011) && ({row_reg, col_reg}<16'b0111100100001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111100100001101) && ({row_reg, col_reg}<16'b0111100100010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111100100010000) && ({row_reg, col_reg}<16'b0111100100010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111100100010100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0111100100010101) && ({row_reg, col_reg}<16'b0111100100011000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111100100011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111100100011001) && ({row_reg, col_reg}<16'b0111100100011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111100100011101) && ({row_reg, col_reg}<16'b0111100100100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111100100100001) && ({row_reg, col_reg}<16'b0111100100100100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111100100100100) && ({row_reg, col_reg}<16'b0111100100100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111100100100110) && ({row_reg, col_reg}<16'b0111100100101001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111100100101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111100100101010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111100100101011) && ({row_reg, col_reg}<16'b0111100100101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111100100101101) && ({row_reg, col_reg}<16'b0111100100101111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111100100101111) && ({row_reg, col_reg}<16'b0111100100110001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111100100110001) && ({row_reg, col_reg}<16'b0111100100111000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111100100111000) && ({row_reg, col_reg}<16'b0111100100111010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111100100111010) && ({row_reg, col_reg}<16'b0111100100111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111100100111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111100100111110) && ({row_reg, col_reg}<16'b0111100101000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111100101000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111100101000001) && ({row_reg, col_reg}<16'b0111100101000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111100101000011) && ({row_reg, col_reg}<16'b0111100101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111100101000110) && ({row_reg, col_reg}<16'b0111100101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111100101001100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111100101001101) && ({row_reg, col_reg}<16'b0111100101011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111100101011000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111100101011001) && ({row_reg, col_reg}<16'b0111100101100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111100101100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111100101100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111100101100010) && ({row_reg, col_reg}<16'b0111100101100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100101100100) && ({row_reg, col_reg}<16'b0111100101100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111100101100110) && ({row_reg, col_reg}<16'b0111100101101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111100101101000) && ({row_reg, col_reg}<16'b0111100101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111100101101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111100101101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111100101101100) && ({row_reg, col_reg}<16'b0111100101101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111100101101110) && ({row_reg, col_reg}<16'b0111100101110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111100101110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111100101110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111100101110011) && ({row_reg, col_reg}<16'b0111100101110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100101110101) && ({row_reg, col_reg}<16'b0111100101110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111100101110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111100101111000) && ({row_reg, col_reg}<16'b0111100101111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100101111100) && ({row_reg, col_reg}<16'b0111100101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111100101111111) && ({row_reg, col_reg}<16'b0111100110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100110000010) && ({row_reg, col_reg}<16'b0111100110000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100110000101) && ({row_reg, col_reg}<16'b0111100110010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100110010011) && ({row_reg, col_reg}<16'b0111100110010110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111100110010110) && ({row_reg, col_reg}<16'b0111100110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111100110011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111100110100000) && ({row_reg, col_reg}<16'b0111100110100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111100110100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111100110100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111100110100100)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==16'b0111100110100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111100110100110) && ({row_reg, col_reg}<16'b0111100110101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111100110101000) && ({row_reg, col_reg}<16'b0111100110110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100110110101) && ({row_reg, col_reg}<16'b0111100110111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111100110111001) && ({row_reg, col_reg}<16'b0111100110111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100110111111) && ({row_reg, col_reg}<16'b0111100111000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111100111000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100111000100) && ({row_reg, col_reg}<16'b0111100111000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111100111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100111001000) && ({row_reg, col_reg}<16'b0111100111001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100111001101) && ({row_reg, col_reg}<16'b0111100111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111100111011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111100111100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100111100001) && ({row_reg, col_reg}<16'b0111100111100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111100111100011) && ({row_reg, col_reg}<16'b0111100111100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100111100101) && ({row_reg, col_reg}<16'b0111100111101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111100111101000) && ({row_reg, col_reg}<16'b0111100111101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100111101011) && ({row_reg, col_reg}<16'b0111100111101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111100111101111) && ({row_reg, col_reg}<16'b0111100111110001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111100111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111100111110010)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0111100111110011) && ({row_reg, col_reg}<16'b0111101000000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101000000000) && ({row_reg, col_reg}<16'b0111101000000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101000000011) && ({row_reg, col_reg}<16'b0111101000000101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111101000000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101000000110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0111101000000111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0111101000001000) && ({row_reg, col_reg}<16'b0111101000001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101000001010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111101000001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111101000001100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111101000001101) && ({row_reg, col_reg}<16'b0111101000010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101000010100) && ({row_reg, col_reg}<16'b0111101000010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111101000010111) && ({row_reg, col_reg}<16'b0111101000011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111101000011010) && ({row_reg, col_reg}<16'b0111101000011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111101000011100) && ({row_reg, col_reg}<16'b0111101000100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101000100000) && ({row_reg, col_reg}<16'b0111101000100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111101000100110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111101000100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111101000101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101000101001) && ({row_reg, col_reg}<16'b0111101000101011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111101000101011) && ({row_reg, col_reg}<16'b0111101000110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101000110001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111101000110010) && ({row_reg, col_reg}<16'b0111101000110100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111101000110100) && ({row_reg, col_reg}<16'b0111101000110111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111101000110111) && ({row_reg, col_reg}<16'b0111101000111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101000111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111101000111100) && ({row_reg, col_reg}<16'b0111101001000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111101001000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111101001000001) && ({row_reg, col_reg}<16'b0111101001001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101001001001) && ({row_reg, col_reg}<16'b0111101001001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111101001001101) && ({row_reg, col_reg}<16'b0111101001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101001010100) && ({row_reg, col_reg}<16'b0111101001011010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111101001011010) && ({row_reg, col_reg}<16'b0111101001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101001011111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111101001100000) && ({row_reg, col_reg}<16'b0111101001100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101001100100) && ({row_reg, col_reg}<16'b0111101001100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111101001100110) && ({row_reg, col_reg}<16'b0111101001101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111101001101010) && ({row_reg, col_reg}<16'b0111101001101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111101001101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111101001101111) && ({row_reg, col_reg}<16'b0111101001110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111101001110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0111101001110011) && ({row_reg, col_reg}<16'b0111101001110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111101001110101) && ({row_reg, col_reg}<16'b0111101001111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111101001111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111101001111001) && ({row_reg, col_reg}<16'b0111101001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111101001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101001111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101001111101) && ({row_reg, col_reg}<16'b0111101010000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101010000011) && ({row_reg, col_reg}<16'b0111101010001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101010001010) && ({row_reg, col_reg}<16'b0111101010010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101010010011) && ({row_reg, col_reg}<16'b0111101010010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101010010101) && ({row_reg, col_reg}<16'b0111101010011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101010011110) && ({row_reg, col_reg}<16'b0111101010100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101010100000) && ({row_reg, col_reg}<16'b0111101010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101010100011) && ({row_reg, col_reg}<16'b0111101010101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101010101101) && ({row_reg, col_reg}<16'b0111101010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101010110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111101010110111) && ({row_reg, col_reg}<16'b0111101010111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101010111001) && ({row_reg, col_reg}<16'b0111101011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101011000000) && ({row_reg, col_reg}<16'b0111101011000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111101011000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101011000100) && ({row_reg, col_reg}<16'b0111101011000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111101011000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101011001000) && ({row_reg, col_reg}<16'b0111101011001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101011001101) && ({row_reg, col_reg}<16'b0111101011010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101011010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101011010011) && ({row_reg, col_reg}<16'b0111101011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101011011111) && ({row_reg, col_reg}<16'b0111101011100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101011100010) && ({row_reg, col_reg}<16'b0111101011100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101011100101) && ({row_reg, col_reg}<16'b0111101011100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111101011100111) && ({row_reg, col_reg}<16'b0111101011101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101011101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101011101011) && ({row_reg, col_reg}<16'b0111101011101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101011101101) && ({row_reg, col_reg}<16'b0111101011110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111101011110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101011110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111101011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111101011110011) && ({row_reg, col_reg}<16'b0111101011110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101011110110) && ({row_reg, col_reg}<16'b0111101011111001)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0111101011111001) && ({row_reg, col_reg}<16'b0111101100000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101100000000) && ({row_reg, col_reg}<16'b0111101100000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101100000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111101100001000) && ({row_reg, col_reg}<16'b0111101100001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101100001011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0111101100001100) && ({row_reg, col_reg}<16'b0111101100001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101100001111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111101100010000) && ({row_reg, col_reg}<16'b0111101100010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101100010100) && ({row_reg, col_reg}<16'b0111101100010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111101100010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101100010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111101100011000) && ({row_reg, col_reg}<16'b0111101100011011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111101100011011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0111101100011100) && ({row_reg, col_reg}<16'b0111101100100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111101100100000) && ({row_reg, col_reg}<16'b0111101100100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101100100010) && ({row_reg, col_reg}<16'b0111101100101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111101100101000) && ({row_reg, col_reg}<16'b0111101100101010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111101100101010) && ({row_reg, col_reg}<16'b0111101100101110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101100101110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111101100101111) && ({row_reg, col_reg}<16'b0111101100110001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111101100110001) && ({row_reg, col_reg}<16'b0111101100110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111101100110011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111101100110100) && ({row_reg, col_reg}<16'b0111101100111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101100111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111101100111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101100111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111101100111011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0111101100111100) && ({row_reg, col_reg}<16'b0111101100111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111101100111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111101101000000) && ({row_reg, col_reg}<16'b0111101101001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101101001000) && ({row_reg, col_reg}<16'b0111101101001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111101101001110) && ({row_reg, col_reg}<16'b0111101101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101101010100) && ({row_reg, col_reg}<16'b0111101101010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111101101010110) && ({row_reg, col_reg}<16'b0111101101011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101101011110) && ({row_reg, col_reg}<16'b0111101101100000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111101101100000) && ({row_reg, col_reg}<16'b0111101101100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101101100010) && ({row_reg, col_reg}<16'b0111101101100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111101101100110) && ({row_reg, col_reg}<16'b0111101101101001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111101101101001) && ({row_reg, col_reg}<16'b0111101101101100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0111101101101100) && ({row_reg, col_reg}<16'b0111101101101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111101101101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111101101110000) && ({row_reg, col_reg}<16'b0111101101110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111101101110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111101101110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111101101110100) && ({row_reg, col_reg}<16'b0111101101110111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0111101101110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111101101111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111101101111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111101101111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101101111011) && ({row_reg, col_reg}<16'b0111101101111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101101111101) && ({row_reg, col_reg}<16'b0111101110000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101110000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111101110000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101110000110) && ({row_reg, col_reg}<16'b0111101110001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101110001001) && ({row_reg, col_reg}<16'b0111101110010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101110010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111101110010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101110010010) && ({row_reg, col_reg}<16'b0111101110010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101110010101) && ({row_reg, col_reg}<16'b0111101110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101110011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101110100000) && ({row_reg, col_reg}<16'b0111101110100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101110100101) && ({row_reg, col_reg}<16'b0111101110101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101110101000) && ({row_reg, col_reg}<16'b0111101110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101110101010) && ({row_reg, col_reg}<16'b0111101110101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101110101101) && ({row_reg, col_reg}<16'b0111101110110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101110110101) && ({row_reg, col_reg}<16'b0111101110111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101110111001) && ({row_reg, col_reg}<16'b0111101110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101110111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111101110111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101111000000) && ({row_reg, col_reg}<16'b0111101111000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111101111000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101111000100) && ({row_reg, col_reg}<16'b0111101111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111101111000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111101111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101111001000) && ({row_reg, col_reg}<16'b0111101111001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101111001101) && ({row_reg, col_reg}<16'b0111101111010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101111010010) && ({row_reg, col_reg}<16'b0111101111010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101111010101) && ({row_reg, col_reg}<16'b0111101111100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101111100101) && ({row_reg, col_reg}<16'b0111101111100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111101111100111) && ({row_reg, col_reg}<16'b0111101111101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101111101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101111101011) && ({row_reg, col_reg}<16'b0111101111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101111110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111101111110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111101111110011) && ({row_reg, col_reg}<16'b0111101111110101)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0111101111110101) && ({row_reg, col_reg}<16'b0111110000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111110000000000) && ({row_reg, col_reg}<16'b0111110000001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110000001001) && ({row_reg, col_reg}<16'b0111110000001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110000001101) && ({row_reg, col_reg}<16'b0111110000001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110000001111) && ({row_reg, col_reg}<16'b0111110000010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111110000010010) && ({row_reg, col_reg}<16'b0111110000011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110000011001) && ({row_reg, col_reg}<16'b0111110000011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110000011101) && ({row_reg, col_reg}<16'b0111110000100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111110000100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110000100010) && ({row_reg, col_reg}<16'b0111110000100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111110000100101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111110000100110) && ({row_reg, col_reg}<16'b0111110000101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111110000101001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111110000101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111110000101011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111110000101100) && ({row_reg, col_reg}<16'b0111110000110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111110000110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111110000110011) && ({row_reg, col_reg}<16'b0111110000110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110000110110) && ({row_reg, col_reg}<16'b0111110000111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110000111110) && ({row_reg, col_reg}<16'b0111110001000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110001000010) && ({row_reg, col_reg}<16'b0111110001000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110001000100) && ({row_reg, col_reg}<16'b0111110001001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110001001001) && ({row_reg, col_reg}<16'b0111110001001111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111110001001111) && ({row_reg, col_reg}<16'b0111110001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110001010100) && ({row_reg, col_reg}<16'b0111110001010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111110001010110) && ({row_reg, col_reg}<16'b0111110001011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111110001011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110001011101) && ({row_reg, col_reg}<16'b0111110001100000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111110001100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110001100001) && ({row_reg, col_reg}<16'b0111110001100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111110001100011) && ({row_reg, col_reg}<16'b0111110001100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110001100101) && ({row_reg, col_reg}<16'b0111110001101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111110001101000) && ({row_reg, col_reg}<16'b0111110001101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111110001101010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0111110001101011) && ({row_reg, col_reg}<16'b0111110001101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110001101101) && ({row_reg, col_reg}<16'b0111110001101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111110001101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110001110000) && ({row_reg, col_reg}<16'b0111110001110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111110001110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0111110001110011) && ({row_reg, col_reg}<16'b0111110001110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111110001110101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0111110001110110) && ({row_reg, col_reg}<16'b0111110001111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111110001111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111110001111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110001111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110001111011) && ({row_reg, col_reg}<16'b0111110010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110010000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110010000010) && ({row_reg, col_reg}<16'b0111110010001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110010001111) && ({row_reg, col_reg}<16'b0111110010010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111110010010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110010010010) && ({row_reg, col_reg}<16'b0111110010011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110010011001) && ({row_reg, col_reg}<16'b0111110010100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110010100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110010100111) && ({row_reg, col_reg}<16'b0111110010110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110010110100) && ({row_reg, col_reg}<16'b0111110010110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111110010110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111110010110111) && ({row_reg, col_reg}<16'b0111110010111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110010111001) && ({row_reg, col_reg}<16'b0111110011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110011000000) && ({row_reg, col_reg}<16'b0111110011000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111110011000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110011000011) && ({row_reg, col_reg}<16'b0111110011000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111110011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111110011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110011000111) && ({row_reg, col_reg}<16'b0111110011001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110011001101) && ({row_reg, col_reg}<16'b0111110011010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110011010011) && ({row_reg, col_reg}<16'b0111110011010110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110011010110) && ({row_reg, col_reg}<16'b0111110011011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110011011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110011011010) && ({row_reg, col_reg}<16'b0111110011100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110011100010) && ({row_reg, col_reg}<16'b0111110011100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111110011100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110011100101) && ({row_reg, col_reg}<16'b0111110011100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111110011100111) && ({row_reg, col_reg}<16'b0111110011101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110011101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110011101110) && ({row_reg, col_reg}<16'b0111110011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110011110001) && ({row_reg, col_reg}<16'b0111110011110100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0111110011110100) && ({row_reg, col_reg}<16'b0111110100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111110100000000) && ({row_reg, col_reg}<16'b0111110100000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111110100000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110100000111) && ({row_reg, col_reg}<16'b0111110100001001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0111110100001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110100001010) && ({row_reg, col_reg}<16'b0111110100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111110100001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111110100001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111110100001111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111110100010000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111110100010001) && ({row_reg, col_reg}<16'b0111110100010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111110100010011) && ({row_reg, col_reg}<16'b0111110100011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110100011001) && ({row_reg, col_reg}<16'b0111110100011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110100011011) && ({row_reg, col_reg}<16'b0111110100011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110100011101) && ({row_reg, col_reg}<16'b0111110100100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111110100100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110100100011) && ({row_reg, col_reg}<16'b0111110100101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111110100101000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111110100101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111110100101010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111110100101011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111110100101100) && ({row_reg, col_reg}<16'b0111110100110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111110100110001) && ({row_reg, col_reg}<16'b0111110100110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111110100110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111110100110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111110100110110) && ({row_reg, col_reg}<16'b0111110100111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111110100111000) && ({row_reg, col_reg}<16'b0111110100111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110100111010) && ({row_reg, col_reg}<16'b0111110101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111110101010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111110101010001) && ({row_reg, col_reg}<16'b0111110101011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110101011001) && ({row_reg, col_reg}<16'b0111110101011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110101011011) && ({row_reg, col_reg}<16'b0111110101011101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111110101011101) && ({row_reg, col_reg}<16'b0111110101100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110101100001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111110101100010) && ({row_reg, col_reg}<16'b0111110101101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110101101100) && ({row_reg, col_reg}<16'b0111110101101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0111110101101111) && ({row_reg, col_reg}<16'b0111110101110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111110101110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0111110101110011) && ({row_reg, col_reg}<16'b0111110101110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111110101110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111110101111000) && ({row_reg, col_reg}<16'b0111110101111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110101111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110101111011) && ({row_reg, col_reg}<16'b0111110110000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110110000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110110001000) && ({row_reg, col_reg}<16'b0111110110001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110110001101) && ({row_reg, col_reg}<16'b0111110110001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110110001111) && ({row_reg, col_reg}<16'b0111110110101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110110101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110110101101) && ({row_reg, col_reg}<16'b0111110110110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110110110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110110110110) && ({row_reg, col_reg}<16'b0111110110111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111110110111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110110111010) && ({row_reg, col_reg}<16'b0111110111000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110111000011) && ({row_reg, col_reg}<16'b0111110111000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111110111000111) && ({row_reg, col_reg}<16'b0111110111001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110111001001) && ({row_reg, col_reg}<16'b0111110111001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110111001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110111001101) && ({row_reg, col_reg}<16'b0111110111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110111010001) && ({row_reg, col_reg}<16'b0111110111010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110111010100) && ({row_reg, col_reg}<16'b0111110111011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110111011000) && ({row_reg, col_reg}<16'b0111110111011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110111011010) && ({row_reg, col_reg}<16'b0111110111011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110111011110) && ({row_reg, col_reg}<16'b0111110111100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110111100000) && ({row_reg, col_reg}<16'b0111110111100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110111100010) && ({row_reg, col_reg}<16'b0111110111100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110111100100) && ({row_reg, col_reg}<16'b0111110111101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110111101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110111101110) && ({row_reg, col_reg}<16'b0111110111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110111110001) && ({row_reg, col_reg}<16'b0111110111110100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0111110111110100) && ({row_reg, col_reg}<16'b0111111000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111111000000000) && ({row_reg, col_reg}<16'b0111111000000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111000000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111000000111) && ({row_reg, col_reg}<16'b0111111000001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111000001010) && ({row_reg, col_reg}<16'b0111111000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111111000001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111000001110) && ({row_reg, col_reg}<16'b0111111000010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111000010000) && ({row_reg, col_reg}<16'b0111111000010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111111000010100) && ({row_reg, col_reg}<16'b0111111000011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111000011101) && ({row_reg, col_reg}<16'b0111111000100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111000100111) && ({row_reg, col_reg}<16'b0111111000101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111000101011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111111000101100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111111000101101) && ({row_reg, col_reg}<16'b0111111000101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111111000101111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111111000110000) && ({row_reg, col_reg}<16'b0111111000110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111000110010) && ({row_reg, col_reg}<16'b0111111000110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111000110101) && ({row_reg, col_reg}<16'b0111111000110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111111000110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111000111000) && ({row_reg, col_reg}<16'b0111111000111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111000111101) && ({row_reg, col_reg}<16'b0111111001000001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111111001000001) && ({row_reg, col_reg}<16'b0111111001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111001010000) && ({row_reg, col_reg}<16'b0111111001010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111111001010010) && ({row_reg, col_reg}<16'b0111111001011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111001011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111001011010) && ({row_reg, col_reg}<16'b0111111001011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111111001011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111001011101) && ({row_reg, col_reg}<16'b0111111001100000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111111001100000) && ({row_reg, col_reg}<16'b0111111001100010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111111001100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111001100011) && ({row_reg, col_reg}<16'b0111111001100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111111001100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111001100110) && ({row_reg, col_reg}<16'b0111111001101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111001101000) && ({row_reg, col_reg}<16'b0111111001101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111111001101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0111111001101011) && ({row_reg, col_reg}<16'b0111111001101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111111001101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0111111001110000) && ({row_reg, col_reg}<16'b0111111001110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111001110010) && ({row_reg, col_reg}<16'b0111111001110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111111001110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111111001110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111111001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111001111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111001111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111001111011) && ({row_reg, col_reg}<16'b0111111001111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111001111101) && ({row_reg, col_reg}<16'b0111111010100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111010100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111111010100110) && ({row_reg, col_reg}<16'b0111111010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111010110110) && ({row_reg, col_reg}<16'b0111111010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111111010111010) && ({row_reg, col_reg}<16'b0111111010111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111111010111110) && ({row_reg, col_reg}<16'b0111111011000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111011000011) && ({row_reg, col_reg}<16'b0111111011000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111111011000111) && ({row_reg, col_reg}<16'b0111111011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111011001010) && ({row_reg, col_reg}<16'b0111111011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111011010001) && ({row_reg, col_reg}<16'b0111111011010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111011010101) && ({row_reg, col_reg}<16'b0111111011011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111011011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111011011010) && ({row_reg, col_reg}<16'b0111111011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111011011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111011100000) && ({row_reg, col_reg}<16'b0111111011100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111011100010) && ({row_reg, col_reg}<16'b0111111011100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111011100100) && ({row_reg, col_reg}<16'b0111111011101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111011101011) && ({row_reg, col_reg}<16'b0111111011101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111011101110) && ({row_reg, col_reg}<16'b0111111011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111011110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111111011110011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0111111011110100) && ({row_reg, col_reg}<16'b0111111100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111111100000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111100000001) && ({row_reg, col_reg}<16'b0111111100000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111100000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111100000110) && ({row_reg, col_reg}<16'b0111111100001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111100001010) && ({row_reg, col_reg}<16'b0111111100001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111100001110) && ({row_reg, col_reg}<16'b0111111100010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111100010000) && ({row_reg, col_reg}<16'b0111111100010101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111111100010101) && ({row_reg, col_reg}<16'b0111111100011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111100011101) && ({row_reg, col_reg}<16'b0111111100011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111100011111) && ({row_reg, col_reg}<16'b0111111100100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111100100011) && ({row_reg, col_reg}<16'b0111111100101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111100101010) && ({row_reg, col_reg}<16'b0111111100110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111100110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111100110010) && ({row_reg, col_reg}<16'b0111111100110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111111100110100) && ({row_reg, col_reg}<16'b0111111100110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111100110111) && ({row_reg, col_reg}<16'b0111111100111100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111100111100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111111100111101) && ({row_reg, col_reg}<16'b0111111101000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111101000000) && ({row_reg, col_reg}<16'b0111111101000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111111101000010) && ({row_reg, col_reg}<16'b0111111101001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111101001111) && ({row_reg, col_reg}<16'b0111111101010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111111101010010) && ({row_reg, col_reg}<16'b0111111101011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111101011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111111101011001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111111101011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111101011011) && ({row_reg, col_reg}<16'b0111111101011111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111111101011111) && ({row_reg, col_reg}<16'b0111111101100001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111111101100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111101100010) && ({row_reg, col_reg}<16'b0111111101100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111111101100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111101100101) && ({row_reg, col_reg}<16'b0111111101101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111101101001) && ({row_reg, col_reg}<16'b0111111101101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111101101110) && ({row_reg, col_reg}<16'b0111111101110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111111101110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111111101110001)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}>=16'b0111111101110010) && ({row_reg, col_reg}<16'b0111111101110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111111101110101)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==16'b0111111101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111111101110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111101111000) && ({row_reg, col_reg}<16'b0111111101111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111101111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111101111011) && ({row_reg, col_reg}<16'b0111111101111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111101111101) && ({row_reg, col_reg}<16'b0111111110001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111110001011) && ({row_reg, col_reg}<16'b0111111110001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111110001101) && ({row_reg, col_reg}<16'b0111111110010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111110010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111110010100) && ({row_reg, col_reg}<16'b0111111110011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111110011011) && ({row_reg, col_reg}<16'b0111111110011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111110011110) && ({row_reg, col_reg}<16'b0111111110110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111110110011) && ({row_reg, col_reg}<16'b0111111110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111111110110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111110110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111111110110111) && ({row_reg, col_reg}<16'b0111111110111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111111110111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111110111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111111000000) && ({row_reg, col_reg}<16'b0111111111000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111111111000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111111000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111111111000100) && ({row_reg, col_reg}<16'b0111111111000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111111111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111111001000) && ({row_reg, col_reg}<16'b0111111111001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111111001010) && ({row_reg, col_reg}<16'b0111111111100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111111100010) && ({row_reg, col_reg}<16'b0111111111100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111111111100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111111100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111111111100110) && ({row_reg, col_reg}<16'b0111111111101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111111101011) && ({row_reg, col_reg}<16'b0111111111101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111111101110) && ({row_reg, col_reg}<16'b0111111111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111111110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111111110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111111111110011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b0111111111110100) && ({row_reg, col_reg}<16'b1000000000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000000000000000) && ({row_reg, col_reg}<16'b1000000000000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000000000011) && ({row_reg, col_reg}<16'b1000000000010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000000010000) && ({row_reg, col_reg}<16'b1000000000010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000000000010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000000010011) && ({row_reg, col_reg}<16'b1000000000010101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000000000010101) && ({row_reg, col_reg}<16'b1000000000100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000000100111) && ({row_reg, col_reg}<16'b1000000000101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000000101101) && ({row_reg, col_reg}<16'b1000000000110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000000000110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000000110010) && ({row_reg, col_reg}<16'b1000000000110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000000000110100) && ({row_reg, col_reg}<16'b1000000000110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000000110110) && ({row_reg, col_reg}<16'b1000000000111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000000111011) && ({row_reg, col_reg}<16'b1000000000111101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000000000111101) && ({row_reg, col_reg}<16'b1000000001001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000001001110) && ({row_reg, col_reg}<16'b1000000001010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000000001010010) && ({row_reg, col_reg}<16'b1000000001010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000000001010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000000001011000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000000001011001) && ({row_reg, col_reg}<16'b1000000001011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000001011011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000000001011100) && ({row_reg, col_reg}<16'b1000000001100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000000001100000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000000001100001) && ({row_reg, col_reg}<16'b1000000001100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000000001100011) && ({row_reg, col_reg}<16'b1000000001100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000001100101) && ({row_reg, col_reg}<16'b1000000001100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000001100111) && ({row_reg, col_reg}<16'b1000000001101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000001101001) && ({row_reg, col_reg}<16'b1000000001101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000000001101100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1000000001101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000000001101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000000001101111) && ({row_reg, col_reg}<16'b1000000001110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000001110010) && ({row_reg, col_reg}<16'b1000000001110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000000001110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000000001110101) && ({row_reg, col_reg}<16'b1000000001110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000000001110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000001111000) && ({row_reg, col_reg}<16'b1000000001111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000000001111010) && ({row_reg, col_reg}<16'b1000000001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000001111100) && ({row_reg, col_reg}<16'b1000000010000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000010000100) && ({row_reg, col_reg}<16'b1000000010000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000010000110) && ({row_reg, col_reg}<16'b1000000010001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000010001000) && ({row_reg, col_reg}<16'b1000000010001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000010001010) && ({row_reg, col_reg}<16'b1000000010010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000010010100) && ({row_reg, col_reg}<16'b1000000010011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000010011001) && ({row_reg, col_reg}<16'b1000000010101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000010101110) && ({row_reg, col_reg}<16'b1000000010110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000010110010) && ({row_reg, col_reg}<16'b1000000010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000000010110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000010110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000000010110111) && ({row_reg, col_reg}<16'b1000000011000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000000011000000) && ({row_reg, col_reg}<16'b1000000011000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000000011000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000011000011) && ({row_reg, col_reg}<16'b1000000011000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000000011000110) && ({row_reg, col_reg}<16'b1000000011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000011001000) && ({row_reg, col_reg}<16'b1000000011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000011001011) && ({row_reg, col_reg}<16'b1000000011100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000011100010) && ({row_reg, col_reg}<16'b1000000011100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000011100100) && ({row_reg, col_reg}<16'b1000000011100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000000011100110) && ({row_reg, col_reg}<16'b1000000011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000011101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000000011110000) && ({row_reg, col_reg}<16'b1000000011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000000011110011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b1000000011110100) && ({row_reg, col_reg}<16'b1000000100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000000100000000) && ({row_reg, col_reg}<16'b1000000100000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000000100000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000100000011) && ({row_reg, col_reg}<16'b1000000100001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000000100001010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000000100001011) && ({row_reg, col_reg}<16'b1000000100010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000000100010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000000100010101) && ({row_reg, col_reg}<16'b1000000100101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000100101000) && ({row_reg, col_reg}<16'b1000000100101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000100101100) && ({row_reg, col_reg}<16'b1000000100101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000000100101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000100101111) && ({row_reg, col_reg}<16'b1000000100110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000100110001) && ({row_reg, col_reg}<16'b1000000100110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000100110111) && ({row_reg, col_reg}<16'b1000000100111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000100111010) && ({row_reg, col_reg}<16'b1000000100111101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000000100111101) && ({row_reg, col_reg}<16'b1000000101001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000101001110) && ({row_reg, col_reg}<16'b1000000101010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000000101010010) && ({row_reg, col_reg}<16'b1000000101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000101010100) && ({row_reg, col_reg}<16'b1000000101010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000101010111) && ({row_reg, col_reg}<16'b1000000101011001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000000101011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000101011010) && ({row_reg, col_reg}<16'b1000000101011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000000101011100) && ({row_reg, col_reg}<16'b1000000101011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000000101011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1000000101100000)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==16'b1000000101100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000000101100010) && ({row_reg, col_reg}<16'b1000000101101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000101101100) && ({row_reg, col_reg}<16'b1000000101101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000000101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000101110000) && ({row_reg, col_reg}<16'b1000000101110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000000101110010) && ({row_reg, col_reg}<16'b1000000101110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000101110100) && ({row_reg, col_reg}<16'b1000000101110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000000101110110) && ({row_reg, col_reg}<16'b1000000101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000101111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000000101111001) && ({row_reg, col_reg}<16'b1000000101111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000101111101) && ({row_reg, col_reg}<16'b1000000110000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000110000100) && ({row_reg, col_reg}<16'b1000000110000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000110000110) && ({row_reg, col_reg}<16'b1000000110001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000110001000) && ({row_reg, col_reg}<16'b1000000110001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000110001010) && ({row_reg, col_reg}<16'b1000000110010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000110010011) && ({row_reg, col_reg}<16'b1000000110010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000110010110) && ({row_reg, col_reg}<16'b1000000110011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000110011110) && ({row_reg, col_reg}<16'b1000000110100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000110100000) && ({row_reg, col_reg}<16'b1000000110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000000110110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000110110110) && ({row_reg, col_reg}<16'b1000000110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000000110111000) && ({row_reg, col_reg}<16'b1000000110111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000000110111011) && ({row_reg, col_reg}<16'b1000000111000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000000111000010) && ({row_reg, col_reg}<16'b1000000111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000000111000110) && ({row_reg, col_reg}<16'b1000000111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000111001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000111001001) && ({row_reg, col_reg}<16'b1000000111100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000111100010) && ({row_reg, col_reg}<16'b1000000111100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000111100100) && ({row_reg, col_reg}<16'b1000000111100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000000111100110) && ({row_reg, col_reg}<16'b1000000111101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000111101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000000111101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000111101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000000111110000) && ({row_reg, col_reg}<16'b1000000111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000111110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000000111110011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b1000000111110100) && ({row_reg, col_reg}<16'b1000001000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000001000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001000000001) && ({row_reg, col_reg}<16'b1000001000000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000001000000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001000000100) && ({row_reg, col_reg}<16'b1000001000001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001000001010) && ({row_reg, col_reg}<16'b1000001000001100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000001000001100) && ({row_reg, col_reg}<16'b1000001000010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001000010000) && ({row_reg, col_reg}<16'b1000001000010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000001000010010) && ({row_reg, col_reg}<16'b1000001000010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000001000010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000001000010101) && ({row_reg, col_reg}<16'b1000001000101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001000101000) && ({row_reg, col_reg}<16'b1000001000101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001000101100) && ({row_reg, col_reg}<16'b1000001000101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000001000101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001000101111) && ({row_reg, col_reg}<16'b1000001000110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001000110001) && ({row_reg, col_reg}<16'b1000001000110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001000110100) && ({row_reg, col_reg}<16'b1000001000111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001000111001) && ({row_reg, col_reg}<16'b1000001000111101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000001000111101) && ({row_reg, col_reg}<16'b1000001001000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001001000100) && ({row_reg, col_reg}<16'b1000001001000110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000001001000110) && ({row_reg, col_reg}<16'b1000001001001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001001001110) && ({row_reg, col_reg}<16'b1000001001010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000001001010010) && ({row_reg, col_reg}<16'b1000001001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001001010100) && ({row_reg, col_reg}<16'b1000001001010111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000001001010111) && ({row_reg, col_reg}<16'b1000001001011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001001011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000001001011011) && ({row_reg, col_reg}<16'b1000001001100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001001100011) && ({row_reg, col_reg}<16'b1000001001100101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1000001001100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000001001100110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000001001100111) && ({row_reg, col_reg}<16'b1000001001101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001001101001) && ({row_reg, col_reg}<16'b1000001001101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1000001001101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000001001101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000001001101101) && ({row_reg, col_reg}<16'b1000001001110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000001001110001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1000001001110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000001001110011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1000001001110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000001001110101) && ({row_reg, col_reg}<16'b1000001001110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001001110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000001001111000) && ({row_reg, col_reg}<16'b1000001001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001001111101) && ({row_reg, col_reg}<16'b1000001010010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001010010011) && ({row_reg, col_reg}<16'b1000001010010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001010010110) && ({row_reg, col_reg}<16'b1000001010011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001010011110) && ({row_reg, col_reg}<16'b1000001010100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001010100001) && ({row_reg, col_reg}<16'b1000001010110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001010110100) && ({row_reg, col_reg}<16'b1000001010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001010110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000001010110111) && ({row_reg, col_reg}<16'b1000001010111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000001010111001) && ({row_reg, col_reg}<16'b1000001010111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001010111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000001010111100) && ({row_reg, col_reg}<16'b1000001011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000001011000011) && ({row_reg, col_reg}<16'b1000001011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001011001000) && ({row_reg, col_reg}<16'b1000001011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001011001010) && ({row_reg, col_reg}<16'b1000001011100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001011100010) && ({row_reg, col_reg}<16'b1000001011100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000001011100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001011100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000001011100110) && ({row_reg, col_reg}<16'b1000001011101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001011101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000001011101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001011101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000001011110000) && ({row_reg, col_reg}<16'b1000001011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000001011110011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b1000001011110100) && ({row_reg, col_reg}<16'b1000001100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000001100000000) && ({row_reg, col_reg}<16'b1000001100000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001100000010) && ({row_reg, col_reg}<16'b1000001100000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000001100000100) && ({row_reg, col_reg}<16'b1000001100001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001100001000) && ({row_reg, col_reg}<16'b1000001100010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000001100010000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000001100010001) && ({row_reg, col_reg}<16'b1000001100010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000001100010110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000001100010111) && ({row_reg, col_reg}<16'b1000001100011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001100011111) && ({row_reg, col_reg}<16'b1000001100100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000001100100001) && ({row_reg, col_reg}<16'b1000001100101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000001100101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001100101010) && ({row_reg, col_reg}<16'b1000001100101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000001100101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000001100101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000001100101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001100101111) && ({row_reg, col_reg}<16'b1000001100110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000001100110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001100110011) && ({row_reg, col_reg}<16'b1000001100111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001100111010) && ({row_reg, col_reg}<16'b1000001100111100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000001100111100) && ({row_reg, col_reg}<16'b1000001101000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000001101000011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000001101000100) && ({row_reg, col_reg}<16'b1000001101000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000001101000110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000001101000111) && ({row_reg, col_reg}<16'b1000001101001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001101001110) && ({row_reg, col_reg}<16'b1000001101010001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000001101010001) && ({row_reg, col_reg}<16'b1000001101010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000001101010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000001101010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000001101010101) && ({row_reg, col_reg}<16'b1000001101011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001101011001) && ({row_reg, col_reg}<16'b1000001101011011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000001101011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000001101011100) && ({row_reg, col_reg}<16'b1000001101100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000001101100110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000001101100111) && ({row_reg, col_reg}<16'b1000001101101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001101101001) && ({row_reg, col_reg}<16'b1000001101101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1000001101101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000001101101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000001101101110) && ({row_reg, col_reg}<16'b1000001101110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000001101110001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1000001101110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000001101110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000001101110100) && ({row_reg, col_reg}<16'b1000001101110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000001101110111) && ({row_reg, col_reg}<16'b1000001101111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001101111001) && ({row_reg, col_reg}<16'b1000001101111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000001101111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001101111101) && ({row_reg, col_reg}<16'b1000001110010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001110010100) && ({row_reg, col_reg}<16'b1000001110011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001110011001) && ({row_reg, col_reg}<16'b1000001110011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001110011011) && ({row_reg, col_reg}<16'b1000001110100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001110100001) && ({row_reg, col_reg}<16'b1000001110110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001110110011) && ({row_reg, col_reg}<16'b1000001110110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001110110110) && ({row_reg, col_reg}<16'b1000001110111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000001110111001) && ({row_reg, col_reg}<16'b1000001110111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001110111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000001110111100)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==16'b1000001110111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000001110111110) && ({row_reg, col_reg}<16'b1000001111000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000001111000000) && ({row_reg, col_reg}<16'b1000001111000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000001111000010)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==16'b1000001111000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001111000100) && ({row_reg, col_reg}<16'b1000001111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001111001001) && ({row_reg, col_reg}<16'b1000001111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001111001011) && ({row_reg, col_reg}<16'b1000001111100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001111100010) && ({row_reg, col_reg}<16'b1000001111100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001111100100) && ({row_reg, col_reg}<16'b1000001111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001111101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000001111110000) && ({row_reg, col_reg}<16'b1000001111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001111110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000001111110011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b1000001111110100) && ({row_reg, col_reg}<16'b1000010000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000010000000000) && ({row_reg, col_reg}<16'b1000010000001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000010000001000) && ({row_reg, col_reg}<16'b1000010000001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010000001010) && ({row_reg, col_reg}<16'b1000010000001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010000001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010000001101) && ({row_reg, col_reg}<16'b1000010000011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000010000011000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010000011001) && ({row_reg, col_reg}<16'b1000010000011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000010000011100) && ({row_reg, col_reg}<16'b1000010000011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010000011110) && ({row_reg, col_reg}<16'b1000010000100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000010000100001) && ({row_reg, col_reg}<16'b1000010000100100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000010000100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000010000100101) && ({row_reg, col_reg}<16'b1000010000100111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010000100111) && ({row_reg, col_reg}<16'b1000010000101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000010000101100) && ({row_reg, col_reg}<16'b1000010000101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010000101110) && ({row_reg, col_reg}<16'b1000010000110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010000110100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000010000110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000010000110110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010000110111) && ({row_reg, col_reg}<16'b1000010000111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000010000111010) && ({row_reg, col_reg}<16'b1000010000111100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000010000111100) && ({row_reg, col_reg}<16'b1000010001000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010001000000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000010001000001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010001000010) && ({row_reg, col_reg}<16'b1000010001000111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000010001000111) && ({row_reg, col_reg}<16'b1000010001001010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010001001010) && ({row_reg, col_reg}<16'b1000010001001100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000010001001100) && ({row_reg, col_reg}<16'b1000010001001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000010001001110) && ({row_reg, col_reg}<16'b1000010001010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000010001010000) && ({row_reg, col_reg}<16'b1000010001010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010001010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000010001010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000010001010100) && ({row_reg, col_reg}<16'b1000010001011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010001011000) && ({row_reg, col_reg}<16'b1000010001011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000010001011010) && ({row_reg, col_reg}<16'b1000010001011101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000010001011101) && ({row_reg, col_reg}<16'b1000010001100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000010001100010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000010001100011) && ({row_reg, col_reg}<16'b1000010001100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000010001100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000010001100110) && ({row_reg, col_reg}<16'b1000010001101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000010001101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1000010001101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010001101011) && ({row_reg, col_reg}<16'b1000010001101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1000010001101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000010001101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000010001101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000010001110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000010001110001) && ({row_reg, col_reg}<16'b1000010001110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000010001110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000010001110100) && ({row_reg, col_reg}<16'b1000010001111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010001111001) && ({row_reg, col_reg}<16'b1000010010001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010010001011) && ({row_reg, col_reg}<16'b1000010010010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010010010000) && ({row_reg, col_reg}<16'b1000010010010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010010010100) && ({row_reg, col_reg}<16'b1000010010011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010010011100) && ({row_reg, col_reg}<16'b1000010010011110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000010010011110) && ({row_reg, col_reg}<16'b1000010010100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010010100001) && ({row_reg, col_reg}<16'b1000010010101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010010101010) && ({row_reg, col_reg}<16'b1000010010101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010010101111) && ({row_reg, col_reg}<16'b1000010010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010010110010) && ({row_reg, col_reg}<16'b1000010010110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010010110111) && ({row_reg, col_reg}<16'b1000010010111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000010010111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010010111011) && ({row_reg, col_reg}<16'b1000010010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010010111101) && ({row_reg, col_reg}<16'b1000010011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010011000000) && ({row_reg, col_reg}<16'b1000010011000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000010011000010) && ({row_reg, col_reg}<16'b1000010011000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010011000110) && ({row_reg, col_reg}<16'b1000010011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010011001001) && ({row_reg, col_reg}<16'b1000010011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010011001011) && ({row_reg, col_reg}<16'b1000010011100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010011100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000010011100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010011100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000010011100110) && ({row_reg, col_reg}<16'b1000010011101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010011101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000010011101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010011101011) && ({row_reg, col_reg}<16'b1000010011101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010011101101) && ({row_reg, col_reg}<16'b1000010011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010011101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000010011110000) && ({row_reg, col_reg}<16'b1000010011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000010011110011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b1000010011110100) && ({row_reg, col_reg}<16'b1000010100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000010100000000) && ({row_reg, col_reg}<16'b1000010100000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000010100000010) && ({row_reg, col_reg}<16'b1000010100001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010100001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000010100001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010100001010) && ({row_reg, col_reg}<16'b1000010100001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010100001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010100001101) && ({row_reg, col_reg}<16'b1000010100010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000010100010010) && ({row_reg, col_reg}<16'b1000010100010101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000010100010101) && ({row_reg, col_reg}<16'b1000010100011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000010100011001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000010100011010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000010100011011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010100011100) && ({row_reg, col_reg}<16'b1000010100101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000010100101000) && ({row_reg, col_reg}<16'b1000010100110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010100110001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000010100110010) && ({row_reg, col_reg}<16'b1000010100110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000010100110111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010100111000) && ({row_reg, col_reg}<16'b1000010100111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000010100111010) && ({row_reg, col_reg}<16'b1000010100111110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000010100111110) && ({row_reg, col_reg}<16'b1000010101000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000010101000001) && ({row_reg, col_reg}<16'b1000010101000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000010101000100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000010101000101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000010101000110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010101000111) && ({row_reg, col_reg}<16'b1000010101001010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000010101001010) && ({row_reg, col_reg}<16'b1000010101001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000010101001110) && ({row_reg, col_reg}<16'b1000010101010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010101010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010101010010) && ({row_reg, col_reg}<16'b1000010101010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000010101010100) && ({row_reg, col_reg}<16'b1000010101010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010101010111) && ({row_reg, col_reg}<16'b1000010101011001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000010101011001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1000010101011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010101011011) && ({row_reg, col_reg}<16'b1000010101011101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000010101011101) && ({row_reg, col_reg}<16'b1000010101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000010101100010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000010101100011) && ({row_reg, col_reg}<16'b1000010101100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010101100111) && ({row_reg, col_reg}<16'b1000010101101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000010101101001) && ({row_reg, col_reg}<16'b1000010101101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000010101101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000010101101101) && ({row_reg, col_reg}<16'b1000010101110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010101110000) && ({row_reg, col_reg}<16'b1000010101110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000010101110010) && ({row_reg, col_reg}<16'b1000010101111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010101111001) && ({row_reg, col_reg}<16'b1000010110000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010110000000) && ({row_reg, col_reg}<16'b1000010110000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010110000011) && ({row_reg, col_reg}<16'b1000010110001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010110001001) && ({row_reg, col_reg}<16'b1000010110011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010110011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010110011001) && ({row_reg, col_reg}<16'b1000010110011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010110011011) && ({row_reg, col_reg}<16'b1000010110011110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000010110011110) && ({row_reg, col_reg}<16'b1000010110100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010110100001) && ({row_reg, col_reg}<16'b1000010110101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010110101010) && ({row_reg, col_reg}<16'b1000010110101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010110101111) && ({row_reg, col_reg}<16'b1000010110110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010110110001) && ({row_reg, col_reg}<16'b1000010110110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010110110111) && ({row_reg, col_reg}<16'b1000010110111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000010110111001) && ({row_reg, col_reg}<16'b1000010110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010110111101) && ({row_reg, col_reg}<16'b1000010110111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000010110111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010111000000) && ({row_reg, col_reg}<16'b1000010111000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000010111000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010111000011) && ({row_reg, col_reg}<16'b1000010111000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010111000110) && ({row_reg, col_reg}<16'b1000010111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010111001000) && ({row_reg, col_reg}<16'b1000010111001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010111001100) && ({row_reg, col_reg}<16'b1000010111011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010111011110) && ({row_reg, col_reg}<16'b1000010111100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010111100000) && ({row_reg, col_reg}<16'b1000010111100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010111100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000010111100110) && ({row_reg, col_reg}<16'b1000010111101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010111101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000010111101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010111101011) && ({row_reg, col_reg}<16'b1000010111101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010111101101) && ({row_reg, col_reg}<16'b1000010111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010111101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000010111110000) && ({row_reg, col_reg}<16'b1000010111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010111110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000010111110011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b1000010111110100) && ({row_reg, col_reg}<16'b1000011000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000011000000000) && ({row_reg, col_reg}<16'b1000011000000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011000000010) && ({row_reg, col_reg}<16'b1000011000001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011000001000) && ({row_reg, col_reg}<16'b1000011000001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000011000001010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000011000001011) && ({row_reg, col_reg}<16'b1000011000001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000011000001101) && ({row_reg, col_reg}<16'b1000011000010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000011000010001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000011000010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000011000010011) && ({row_reg, col_reg}<16'b1000011000010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000011000010101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000011000010110) && ({row_reg, col_reg}<16'b1000011000011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000011000011001) && ({row_reg, col_reg}<16'b1000011000011011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000011000011011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000011000011100) && ({row_reg, col_reg}<16'b1000011000101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000011000101000) && ({row_reg, col_reg}<16'b1000011000101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000011000101111) && ({row_reg, col_reg}<16'b1000011000110001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000011000110001) && ({row_reg, col_reg}<16'b1000011000110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000011000110111) && ({row_reg, col_reg}<16'b1000011000111001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000011000111001) && ({row_reg, col_reg}<16'b1000011000111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000011000111011) && ({row_reg, col_reg}<16'b1000011000111110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000011000111110) && ({row_reg, col_reg}<16'b1000011001000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000011001000001) && ({row_reg, col_reg}<16'b1000011001000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000011001000100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000011001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000011001000110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000011001000111) && ({row_reg, col_reg}<16'b1000011001001010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000011001001010) && ({row_reg, col_reg}<16'b1000011001001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000011001001101) && ({row_reg, col_reg}<16'b1000011001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000011001010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000011001010001) && ({row_reg, col_reg}<16'b1000011001010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011001010100) && ({row_reg, col_reg}<16'b1000011001010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000011001010111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000011001011000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000011001011001) && ({row_reg, col_reg}<16'b1000011001011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000011001011100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000011001011101)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==16'b1000011001011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000011001011111) && ({row_reg, col_reg}<16'b1000011001100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000011001100001) && ({row_reg, col_reg}<16'b1000011001100011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000011001100011) && ({row_reg, col_reg}<16'b1000011001101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000011001101010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000011001101011) && ({row_reg, col_reg}<16'b1000011001110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000011001110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000011001110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000011001110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000011001110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000011001110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011001110101) && ({row_reg, col_reg}<16'b1000011001110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011001110111) && ({row_reg, col_reg}<16'b1000011001111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011001111001) && ({row_reg, col_reg}<16'b1000011001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011001111011) && ({row_reg, col_reg}<16'b1000011001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011001111101) && ({row_reg, col_reg}<16'b1000011001111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011001111111) && ({row_reg, col_reg}<16'b1000011010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011010000001) && ({row_reg, col_reg}<16'b1000011010000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000011010000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011010000100) && ({row_reg, col_reg}<16'b1000011010001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011010001010) && ({row_reg, col_reg}<16'b1000011010010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011010010011) && ({row_reg, col_reg}<16'b1000011010010110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011010010110) && ({row_reg, col_reg}<16'b1000011010011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011010011011) && ({row_reg, col_reg}<16'b1000011010011101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011010011101) && ({row_reg, col_reg}<16'b1000011010100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011010100001) && ({row_reg, col_reg}<16'b1000011010100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011010100110) && ({row_reg, col_reg}<16'b1000011010101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000011010101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000011010101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011010101010) && ({row_reg, col_reg}<16'b1000011010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000011010101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011010101110) && ({row_reg, col_reg}<16'b1000011010110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011010110011) && ({row_reg, col_reg}<16'b1000011010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011010110101) && ({row_reg, col_reg}<16'b1000011010110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011010110111) && ({row_reg, col_reg}<16'b1000011010111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000011010111001) && ({row_reg, col_reg}<16'b1000011010111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011010111100) && ({row_reg, col_reg}<16'b1000011011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011011000000) && ({row_reg, col_reg}<16'b1000011011000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000011011000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000011011000011) && ({row_reg, col_reg}<16'b1000011011000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011011000101) && ({row_reg, col_reg}<16'b1000011011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011011001000) && ({row_reg, col_reg}<16'b1000011011001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011011001101) && ({row_reg, col_reg}<16'b1000011011010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011011010010) && ({row_reg, col_reg}<16'b1000011011010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000011011010101) && ({row_reg, col_reg}<16'b1000011011011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011011011110) && ({row_reg, col_reg}<16'b1000011011100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011011100000) && ({row_reg, col_reg}<16'b1000011011100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000011011100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011011100110) && ({row_reg, col_reg}<16'b1000011011101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011011101011) && ({row_reg, col_reg}<16'b1000011011101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011011101101) && ({row_reg, col_reg}<16'b1000011011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000011011101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011011110000) && ({row_reg, col_reg}<16'b1000011011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000011011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000011011110011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b1000011011110100) && ({row_reg, col_reg}<16'b1000011100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000011100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000011100000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000011100000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011100000011) && ({row_reg, col_reg}<16'b1000011100001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011100001001) && ({row_reg, col_reg}<16'b1000011100001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000011100001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000011100001101) && ({row_reg, col_reg}<16'b1000011100010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000011100010001) && ({row_reg, col_reg}<16'b1000011100011111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000011100011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000011100100000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000011100100001) && ({row_reg, col_reg}<16'b1000011100100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000011100100011) && ({row_reg, col_reg}<16'b1000011100101000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000011100101000) && ({row_reg, col_reg}<16'b1000011100101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000011100101101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000011100101110) && ({row_reg, col_reg}<16'b1000011100110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000011100110101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000011100110110) && ({row_reg, col_reg}<16'b1000011100111000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000011100111000) && ({row_reg, col_reg}<16'b1000011101000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000011101000000) && ({row_reg, col_reg}<16'b1000011101000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000011101000010) && ({row_reg, col_reg}<16'b1000011101000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000011101000100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000011101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000011101000110) && ({row_reg, col_reg}<16'b1000011101001100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000011101001100) && ({row_reg, col_reg}<16'b1000011101001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000011101001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000011101001111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000011101010000) && ({row_reg, col_reg}<16'b1000011101010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011101010010) && ({row_reg, col_reg}<16'b1000011101010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011101010110) && ({row_reg, col_reg}<16'b1000011101011000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000011101011000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000011101011001) && ({row_reg, col_reg}<16'b1000011101011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000011101011100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000011101011101) && ({row_reg, col_reg}<16'b1000011101011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011101011111) && ({row_reg, col_reg}<16'b1000011101100001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000011101100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011101100010) && ({row_reg, col_reg}<16'b1000011101100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000011101100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011101100110) && ({row_reg, col_reg}<16'b1000011101110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000011101110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000011101110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011101110010) && ({row_reg, col_reg}<16'b1000011101110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000011101110100) && ({row_reg, col_reg}<16'b1000011101110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011101110110) && ({row_reg, col_reg}<16'b1000011101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011101111011) && ({row_reg, col_reg}<16'b1000011101111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000011101111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011101111110) && ({row_reg, col_reg}<16'b1000011110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011110000001) && ({row_reg, col_reg}<16'b1000011110000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000011110000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011110000101) && ({row_reg, col_reg}<16'b1000011110001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011110001111) && ({row_reg, col_reg}<16'b1000011110010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011110010011) && ({row_reg, col_reg}<16'b1000011110010110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011110010110) && ({row_reg, col_reg}<16'b1000011110011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011110011101) && ({row_reg, col_reg}<16'b1000011110100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011110100110) && ({row_reg, col_reg}<16'b1000011110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011110101001) && ({row_reg, col_reg}<16'b1000011110101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011110101111) && ({row_reg, col_reg}<16'b1000011110110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011110110010) && ({row_reg, col_reg}<16'b1000011110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000011110110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000011110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000011110110111) && ({row_reg, col_reg}<16'b1000011110111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000011110111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011110111011) && ({row_reg, col_reg}<16'b1000011111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011111000000) && ({row_reg, col_reg}<16'b1000011111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000011111000011) && ({row_reg, col_reg}<16'b1000011111000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011111000110) && ({row_reg, col_reg}<16'b1000011111001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011111001101) && ({row_reg, col_reg}<16'b1000011111010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011111010011) && ({row_reg, col_reg}<16'b1000011111010110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000011111010110) && ({row_reg, col_reg}<16'b1000011111011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011111011110) && ({row_reg, col_reg}<16'b1000011111100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011111100000) && ({row_reg, col_reg}<16'b1000011111100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011111100010) && ({row_reg, col_reg}<16'b1000011111100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011111100100) && ({row_reg, col_reg}<16'b1000011111101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011111101010) && ({row_reg, col_reg}<16'b1000011111101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011111101101) && ({row_reg, col_reg}<16'b1000011111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000011111101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011111110000) && ({row_reg, col_reg}<16'b1000011111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000011111110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000011111110011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b1000011111110100) && ({row_reg, col_reg}<16'b1000100000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000100000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000100000000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000100000000010) && ({row_reg, col_reg}<16'b1000100000010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000100000010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000100000010001) && ({row_reg, col_reg}<16'b1000100000010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000100000010100) && ({row_reg, col_reg}<16'b1000100000010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000100000010110) && ({row_reg, col_reg}<16'b1000100000011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000100000011010) && ({row_reg, col_reg}<16'b1000100000011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000100000011100) && ({row_reg, col_reg}<16'b1000100000011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100000011111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000100000100000) && ({row_reg, col_reg}<16'b1000100000100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000100000100011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000100000100100) && ({row_reg, col_reg}<16'b1000100000100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100000100110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000100000100111) && ({row_reg, col_reg}<16'b1000100000101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000100000101101) && ({row_reg, col_reg}<16'b1000100000110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000100000110110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000100000110111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000100000111000) && ({row_reg, col_reg}<16'b1000100000111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100000111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000100001000000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000100001000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100001000010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000100001000011) && ({row_reg, col_reg}<16'b1000100001000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000100001000101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000100001000110) && ({row_reg, col_reg}<16'b1000100001001001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000100001001001) && ({row_reg, col_reg}<16'b1000100001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100001001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000100001001101) && ({row_reg, col_reg}<16'b1000100001010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000100001010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000100001010101) && ({row_reg, col_reg}<16'b1000100001011001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000100001011001) && ({row_reg, col_reg}<16'b1000100001011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000100001011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000100001011100) && ({row_reg, col_reg}<16'b1000100001100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000100001100000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000100001100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000100001100010) && ({row_reg, col_reg}<16'b1000100001100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100001100101) && ({row_reg, col_reg}<16'b1000100001100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000100001100111) && ({row_reg, col_reg}<16'b1000100001101010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000100001101010) && ({row_reg, col_reg}<16'b1000100001101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000100001101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000100001101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000100001101110) && ({row_reg, col_reg}<16'b1000100001110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000100001110000) && ({row_reg, col_reg}<16'b1000100001110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100001110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100001110011) && ({row_reg, col_reg}<16'b1000100001110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100001110101) && ({row_reg, col_reg}<16'b1000100001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100001111011) && ({row_reg, col_reg}<16'b1000100001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100001111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100001111110) && ({row_reg, col_reg}<16'b1000100010001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100010001100) && ({row_reg, col_reg}<16'b1000100010001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100010001111) && ({row_reg, col_reg}<16'b1000100010011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100010011100) && ({row_reg, col_reg}<16'b1000100010100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100010100110) && ({row_reg, col_reg}<16'b1000100010110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100010110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000100010110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000100010110111) && ({row_reg, col_reg}<16'b1000100010111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100010111010) && ({row_reg, col_reg}<16'b1000100010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100010111110) && ({row_reg, col_reg}<16'b1000100011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100011000000) && ({row_reg, col_reg}<16'b1000100011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000100011000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100011000100) && ({row_reg, col_reg}<16'b1000100011000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100011000111) && ({row_reg, col_reg}<16'b1000100011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000100011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100011001011) && ({row_reg, col_reg}<16'b1000100011001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100011001101) && ({row_reg, col_reg}<16'b1000100011010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100011010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000100011010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100011010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100011010101) && ({row_reg, col_reg}<16'b1000100011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100011011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100011100000) && ({row_reg, col_reg}<16'b1000100011100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100011100010) && ({row_reg, col_reg}<16'b1000100011100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100011100100) && ({row_reg, col_reg}<16'b1000100011101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100011101010) && ({row_reg, col_reg}<16'b1000100011101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100011101101) && ({row_reg, col_reg}<16'b1000100011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100011101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000100011110000) && ({row_reg, col_reg}<16'b1000100011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000100011110011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b1000100011110100) && ({row_reg, col_reg}<16'b1000100100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000100100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000100100000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000100100000010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000100100000011) && ({row_reg, col_reg}<16'b1000100100000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000100100000111) && ({row_reg, col_reg}<16'b1000100100001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000100100001010) && ({row_reg, col_reg}<16'b1000100100001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000100100001101) && ({row_reg, col_reg}<16'b1000100100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100100001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000100100010000) && ({row_reg, col_reg}<16'b1000100100010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000100100010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100100010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000100100010101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000100100010110) && ({row_reg, col_reg}<16'b1000100100011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000100100011010) && ({row_reg, col_reg}<16'b1000100100011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000100100011100) && ({row_reg, col_reg}<16'b1000100100011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100100011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000100100011111) && ({row_reg, col_reg}<16'b1000100100100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000100100100011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000100100100100) && ({row_reg, col_reg}<16'b1000100100100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000100100100110) && ({row_reg, col_reg}<16'b1000100100101000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000100100101000) && ({row_reg, col_reg}<16'b1000100100101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100100101101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000100100101110) && ({row_reg, col_reg}<16'b1000100100110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000100100110111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000100100111000) && ({row_reg, col_reg}<16'b1000100100111100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000100100111100) && ({row_reg, col_reg}<16'b1000100100111110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000100100111110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000100100111111) && ({row_reg, col_reg}<16'b1000100101000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000100101000001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000100101000010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000100101000011) && ({row_reg, col_reg}<16'b1000100101000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000100101000110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000100101000111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000100101001000) && ({row_reg, col_reg}<16'b1000100101001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000100101001100) && ({row_reg, col_reg}<16'b1000100101001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000100101001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100101001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000100101010000) && ({row_reg, col_reg}<16'b1000100101010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000100101010011) && ({row_reg, col_reg}<16'b1000100101010101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000100101010101) && ({row_reg, col_reg}<16'b1000100101010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000100101010111) && ({row_reg, col_reg}<16'b1000100101011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000100101011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100101011101) && ({row_reg, col_reg}<16'b1000100101100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100101100101) && ({row_reg, col_reg}<16'b1000100101101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000100101101000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000100101101001) && ({row_reg, col_reg}<16'b1000100101101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000100101101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000100101101100) && ({row_reg, col_reg}<16'b1000100101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100101101111) && ({row_reg, col_reg}<16'b1000100101110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100101110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100101110010) && ({row_reg, col_reg}<16'b1000100101110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100101110100) && ({row_reg, col_reg}<16'b1000100101111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100101111110) && ({row_reg, col_reg}<16'b1000100110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100110000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100110000010) && ({row_reg, col_reg}<16'b1000100110001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100110001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100110001011) && ({row_reg, col_reg}<16'b1000100110001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100110001101) && ({row_reg, col_reg}<16'b1000100110001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000100110001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100110010000) && ({row_reg, col_reg}<16'b1000100110010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000100110010010) && ({row_reg, col_reg}<16'b1000100110010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100110010100) && ({row_reg, col_reg}<16'b1000100110011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100110011000) && ({row_reg, col_reg}<16'b1000100110011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100110011011) && ({row_reg, col_reg}<16'b1000100110101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100110101001) && ({row_reg, col_reg}<16'b1000100110110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100110110101) && ({row_reg, col_reg}<16'b1000100110111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100110111001) && ({row_reg, col_reg}<16'b1000100110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100110111110) && ({row_reg, col_reg}<16'b1000100111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100111000000) && ({row_reg, col_reg}<16'b1000100111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000100111000011) && ({row_reg, col_reg}<16'b1000100111000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100111000101) && ({row_reg, col_reg}<16'b1000100111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100111001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100111001001) && ({row_reg, col_reg}<16'b1000100111001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100111001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100111001101) && ({row_reg, col_reg}<16'b1000100111010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100111010010) && ({row_reg, col_reg}<16'b1000100111010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100111010101) && ({row_reg, col_reg}<16'b1000100111011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100111011110) && ({row_reg, col_reg}<16'b1000100111100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100111100000) && ({row_reg, col_reg}<16'b1000100111100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100111100010) && ({row_reg, col_reg}<16'b1000100111100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100111100100) && ({row_reg, col_reg}<16'b1000100111101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100111101010) && ({row_reg, col_reg}<16'b1000100111101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100111101101) && ({row_reg, col_reg}<16'b1000100111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100111101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000100111110000) && ({row_reg, col_reg}<16'b1000100111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100111110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000100111110011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b1000100111110100) && ({row_reg, col_reg}<16'b1000101000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000101000000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000101000000001) && ({row_reg, col_reg}<16'b1000101000000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101000000100) && ({row_reg, col_reg}<16'b1000101000000111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000101000000111) && ({row_reg, col_reg}<16'b1000101000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000101000001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000101000001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101000001011) && ({row_reg, col_reg}<16'b1000101000001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000101000001101) && ({row_reg, col_reg}<16'b1000101000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101000010000) && ({row_reg, col_reg}<16'b1000101000010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000101000010011) && ({row_reg, col_reg}<16'b1000101000010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000101000010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101000011000) && ({row_reg, col_reg}<16'b1000101000011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000101000011011) && ({row_reg, col_reg}<16'b1000101000011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000101000011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000101000011111) && ({row_reg, col_reg}<16'b1000101000100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000101000100011) && ({row_reg, col_reg}<16'b1000101000100101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000101000100101) && ({row_reg, col_reg}<16'b1000101000100111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000101000100111) && ({row_reg, col_reg}<16'b1000101000101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000101000101101) && ({row_reg, col_reg}<16'b1000101000101111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000101000101111) && ({row_reg, col_reg}<16'b1000101000110010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000101000110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000101000110011) && ({row_reg, col_reg}<16'b1000101000110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000101000110101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000101000110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000101000110111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000101000111000) && ({row_reg, col_reg}<16'b1000101000111100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000101000111100) && ({row_reg, col_reg}<16'b1000101000111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000101000111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000101001000000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000101001000001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000101001000010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000101001000011) && ({row_reg, col_reg}<16'b1000101001000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000101001000110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000101001000111) && ({row_reg, col_reg}<16'b1000101001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000101001001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101001001011) && ({row_reg, col_reg}<16'b1000101001001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000101001001101) && ({row_reg, col_reg}<16'b1000101001001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000101001001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000101001010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000101001010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000101001010010) && ({row_reg, col_reg}<16'b1000101001011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000101001011000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000101001011001) && ({row_reg, col_reg}<16'b1000101001011100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000101001011100) && ({row_reg, col_reg}<16'b1000101001100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101001100010) && ({row_reg, col_reg}<16'b1000101001101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000101001101000) && ({row_reg, col_reg}<16'b1000101001101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000101001101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000101001101011) && ({row_reg, col_reg}<16'b1000101001101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101001101110) && ({row_reg, col_reg}<16'b1000101001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101001110000) && ({row_reg, col_reg}<16'b1000101001110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101001110010) && ({row_reg, col_reg}<16'b1000101001110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101001110100) && ({row_reg, col_reg}<16'b1000101001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000101001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101001111100) && ({row_reg, col_reg}<16'b1000101001111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101001111110) && ({row_reg, col_reg}<16'b1000101010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101010000001) && ({row_reg, col_reg}<16'b1000101010000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101010000011) && ({row_reg, col_reg}<16'b1000101010001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101010001001) && ({row_reg, col_reg}<16'b1000101010001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101010001100) && ({row_reg, col_reg}<16'b1000101010011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101010011110) && ({row_reg, col_reg}<16'b1000101010101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101010101001) && ({row_reg, col_reg}<16'b1000101010110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101010110101) && ({row_reg, col_reg}<16'b1000101010111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101010111001) && ({row_reg, col_reg}<16'b1000101010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101010111110) && ({row_reg, col_reg}<16'b1000101011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101011000000) && ({row_reg, col_reg}<16'b1000101011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000101011000011) && ({row_reg, col_reg}<16'b1000101011000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101011000101) && ({row_reg, col_reg}<16'b1000101011010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000101011010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000101011010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101011010100) && ({row_reg, col_reg}<16'b1000101011010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101011010110) && ({row_reg, col_reg}<16'b1000101011011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101011011101) && ({row_reg, col_reg}<16'b1000101011100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101011100000) && ({row_reg, col_reg}<16'b1000101011101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101011101010) && ({row_reg, col_reg}<16'b1000101011101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101011101110) && ({row_reg, col_reg}<16'b1000101011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101011110001) && ({row_reg, col_reg}<16'b1000101011110100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b1000101011110100) && ({row_reg, col_reg}<16'b1000101100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000101100000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000101100000001) && ({row_reg, col_reg}<16'b1000101100000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101100000011) && ({row_reg, col_reg}<16'b1000101100000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000101100000101) && ({row_reg, col_reg}<16'b1000101100001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000101100001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000101100001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000101100001010) && ({row_reg, col_reg}<16'b1000101100001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101100001101) && ({row_reg, col_reg}<16'b1000101100001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000101100001111) && ({row_reg, col_reg}<16'b1000101100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101100010001) && ({row_reg, col_reg}<16'b1000101100010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000101100010011) && ({row_reg, col_reg}<16'b1000101100011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101100011000) && ({row_reg, col_reg}<16'b1000101100011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000101100011011) && ({row_reg, col_reg}<16'b1000101100011111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000101100011111) && ({row_reg, col_reg}<16'b1000101100100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000101100100010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000101100100011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000101100100100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000101100100101) && ({row_reg, col_reg}<16'b1000101100100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000101100100111) && ({row_reg, col_reg}<16'b1000101100101010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000101100101010) && ({row_reg, col_reg}<16'b1000101100101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000101100101101) && ({row_reg, col_reg}<16'b1000101100110001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000101100110001) && ({row_reg, col_reg}<16'b1000101100110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000101100110110) && ({row_reg, col_reg}<16'b1000101100111110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000101100111110) && ({row_reg, col_reg}<16'b1000101101000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000101101000010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000101101000011) && ({row_reg, col_reg}<16'b1000101101000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000101101000110) && ({row_reg, col_reg}<16'b1000101101001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000101101001000) && ({row_reg, col_reg}<16'b1000101101001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101101001010) && ({row_reg, col_reg}<16'b1000101101001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000101101001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000101101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000101101010001) && ({row_reg, col_reg}<16'b1000101101010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000101101010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000101101010100) && ({row_reg, col_reg}<16'b1000101101010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000101101010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000101101011000) && ({row_reg, col_reg}<16'b1000101101011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000101101011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000101101011100) && ({row_reg, col_reg}<16'b1000101101100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000101101100001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000101101100010) && ({row_reg, col_reg}<16'b1000101101100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000101101100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000101101100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000101101100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000101101101000) && ({row_reg, col_reg}<16'b1000101101101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000101101101100) && ({row_reg, col_reg}<16'b1000101101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101101101110) && ({row_reg, col_reg}<16'b1000101101110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000101101110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101101110010) && ({row_reg, col_reg}<16'b1000101101110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101101110100) && ({row_reg, col_reg}<16'b1000101101111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101101111010) && ({row_reg, col_reg}<16'b1000101101111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000101101111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101101111110) && ({row_reg, col_reg}<16'b1000101110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101110000001) && ({row_reg, col_reg}<16'b1000101110000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101110000100) && ({row_reg, col_reg}<16'b1000101110000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101110000110) && ({row_reg, col_reg}<16'b1000101110001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101110001000) && ({row_reg, col_reg}<16'b1000101110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101110011111) && ({row_reg, col_reg}<16'b1000101110101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101110101001) && ({row_reg, col_reg}<16'b1000101110101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000101110101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101110101101) && ({row_reg, col_reg}<16'b1000101110110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101110110000) && ({row_reg, col_reg}<16'b1000101110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000101110110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000101110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000101110110111) && ({row_reg, col_reg}<16'b1000101110111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101110111001) && ({row_reg, col_reg}<16'b1000101110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101110111101) && ({row_reg, col_reg}<16'b1000101111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101111000000) && ({row_reg, col_reg}<16'b1000101111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000101111000011) && ({row_reg, col_reg}<16'b1000101111000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101111000101) && ({row_reg, col_reg}<16'b1000101111001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000101111001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101111001011) && ({row_reg, col_reg}<16'b1000101111010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101111010101) && ({row_reg, col_reg}<16'b1000101111010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101111010111) && ({row_reg, col_reg}<16'b1000101111011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101111011101) && ({row_reg, col_reg}<16'b1000101111100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101111100000) && ({row_reg, col_reg}<16'b1000101111101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101111101010) && ({row_reg, col_reg}<16'b1000101111101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101111101111) && ({row_reg, col_reg}<16'b1000101111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101111110001) && ({row_reg, col_reg}<16'b1000101111110100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b1000101111110100) && ({row_reg, col_reg}<16'b1000110000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000110000000000) && ({row_reg, col_reg}<16'b1000110000000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110000000011) && ({row_reg, col_reg}<16'b1000110000000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1000110000000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110000000110) && ({row_reg, col_reg}<16'b1000110000001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000110000001000) && ({row_reg, col_reg}<16'b1000110000001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000110000001101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000110000001110) && ({row_reg, col_reg}<16'b1000110000010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000110000010000) && ({row_reg, col_reg}<16'b1000110000010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110000010011) && ({row_reg, col_reg}<16'b1000110000011000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000110000011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110000011001) && ({row_reg, col_reg}<16'b1000110000011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110000011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000110000011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110000011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110000011111) && ({row_reg, col_reg}<16'b1000110000100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000110000100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000110000100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110000100100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000110000100101) && ({row_reg, col_reg}<16'b1000110000100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000110000100111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000110000101000) && ({row_reg, col_reg}<16'b1000110000101010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000110000101010) && ({row_reg, col_reg}<16'b1000110000101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110000101101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110000101110) && ({row_reg, col_reg}<16'b1000110000110000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000110000110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110000110001) && ({row_reg, col_reg}<16'b1000110000110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000110000110100) && ({row_reg, col_reg}<16'b1000110000110110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000110000110110) && ({row_reg, col_reg}<16'b1000110000111011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000110000111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000110000111100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000110000111101) && ({row_reg, col_reg}<16'b1000110001000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110001000001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000110001000010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000110001000011) && ({row_reg, col_reg}<16'b1000110001000101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000110001000101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000110001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110001000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000110001001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000110001001001) && ({row_reg, col_reg}<16'b1000110001001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110001001011) && ({row_reg, col_reg}<16'b1000110001001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000110001001111) && ({row_reg, col_reg}<16'b1000110001010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110001010010) && ({row_reg, col_reg}<16'b1000110001010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000110001010100) && ({row_reg, col_reg}<16'b1000110001010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110001010110) && ({row_reg, col_reg}<16'b1000110001011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000110001011001) && ({row_reg, col_reg}<16'b1000110001011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110001011011) && ({row_reg, col_reg}<16'b1000110001011111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000110001011111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000110001100000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000110001100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110001100010) && ({row_reg, col_reg}<16'b1000110001100100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000110001100100) && ({row_reg, col_reg}<16'b1000110001100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000110001100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1000110001100111)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b1000110001101000) && ({row_reg, col_reg}<16'b1000110001101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000110001101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110001101101) && ({row_reg, col_reg}<16'b1000110001101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110001101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000110001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110001110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000110001110010) && ({row_reg, col_reg}<16'b1000110001110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110001110100) && ({row_reg, col_reg}<16'b1000110001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110001111011) && ({row_reg, col_reg}<16'b1000110001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110001111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110001111110) && ({row_reg, col_reg}<16'b1000110010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110010000000) && ({row_reg, col_reg}<16'b1000110010000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110010000100) && ({row_reg, col_reg}<16'b1000110010000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110010000110) && ({row_reg, col_reg}<16'b1000110010001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110010001001) && ({row_reg, col_reg}<16'b1000110010100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110010100000) && ({row_reg, col_reg}<16'b1000110010101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110010101001) && ({row_reg, col_reg}<16'b1000110010101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110010101100) && ({row_reg, col_reg}<16'b1000110010101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000110010101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110010101111) && ({row_reg, col_reg}<16'b1000110010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000110010110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110010110011) && ({row_reg, col_reg}<16'b1000110010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000110010110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000110010110111) && ({row_reg, col_reg}<16'b1000110010111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000110010111001) && ({row_reg, col_reg}<16'b1000110010111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110010111101) && ({row_reg, col_reg}<16'b1000110011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110011000000) && ({row_reg, col_reg}<16'b1000110011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000110011000011) && ({row_reg, col_reg}<16'b1000110011000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000110011000101) && ({row_reg, col_reg}<16'b1000110011000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110011000111) && ({row_reg, col_reg}<16'b1000110011001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000110011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110011001011) && ({row_reg, col_reg}<16'b1000110011001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110011001111) && ({row_reg, col_reg}<16'b1000110011010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110011010001) && ({row_reg, col_reg}<16'b1000110011010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110011010101) && ({row_reg, col_reg}<16'b1000110011010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110011010111) && ({row_reg, col_reg}<16'b1000110011011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110011011101) && ({row_reg, col_reg}<16'b1000110011011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000110011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110011100000) && ({row_reg, col_reg}<16'b1000110011100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000110011100010) && ({row_reg, col_reg}<16'b1000110011101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110011101010) && ({row_reg, col_reg}<16'b1000110011101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110011101110) && ({row_reg, col_reg}<16'b1000110011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110011110001) && ({row_reg, col_reg}<16'b1000110011110100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b1000110011110100) && ({row_reg, col_reg}<16'b1000110100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000110100000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000110100000001) && ({row_reg, col_reg}<16'b1000110100000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110100000101) && ({row_reg, col_reg}<16'b1000110100001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000110100001010) && ({row_reg, col_reg}<16'b1000110100001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000110100001110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000110100001111) && ({row_reg, col_reg}<16'b1000110100010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000110100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110100010010) && ({row_reg, col_reg}<16'b1000110100010111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000110100010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110100011000) && ({row_reg, col_reg}<16'b1000110100011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000110100011010) && ({row_reg, col_reg}<16'b1000110100011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000110100011111) && ({row_reg, col_reg}<16'b1000110100100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000110100100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000110100100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110100100011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000110100100100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000110100100101) && ({row_reg, col_reg}<16'b1000110100101010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000110100101010) && ({row_reg, col_reg}<16'b1000110100101110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000110100101110) && ({row_reg, col_reg}<16'b1000110100110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000110100110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110100110001) && ({row_reg, col_reg}<16'b1000110100110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110100110011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000110100110100) && ({row_reg, col_reg}<16'b1000110100110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000110100110110) && ({row_reg, col_reg}<16'b1000110100111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110100111010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110100111011) && ({row_reg, col_reg}<16'b1000110100111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000110100111101) && ({row_reg, col_reg}<16'b1000110101000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000110101000001) && ({row_reg, col_reg}<16'b1000110101000011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110101000011) && ({row_reg, col_reg}<16'b1000110101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000110101000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000110101001000) && ({row_reg, col_reg}<16'b1000110101001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110101001011) && ({row_reg, col_reg}<16'b1000110101001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000110101001101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000110101001110) && ({row_reg, col_reg}<16'b1000110101011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110101011011) && ({row_reg, col_reg}<16'b1000110101011101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000110101011101) && ({row_reg, col_reg}<16'b1000110101100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110101100101) && ({row_reg, col_reg}<16'b1000110101101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1000110101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000110101101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000110101101100) && ({row_reg, col_reg}<16'b1000110101101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110101101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000110101110000) && ({row_reg, col_reg}<16'b1000110101110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110101110100) && ({row_reg, col_reg}<16'b1000110110000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110110000100) && ({row_reg, col_reg}<16'b1000110110000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110110000111) && ({row_reg, col_reg}<16'b1000110110001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110110001011) && ({row_reg, col_reg}<16'b1000110110001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110110001110) && ({row_reg, col_reg}<16'b1000110110011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110110011100) && ({row_reg, col_reg}<16'b1000110110100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110110100000) && ({row_reg, col_reg}<16'b1000110110101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110110101001) && ({row_reg, col_reg}<16'b1000110110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110110101101) && ({row_reg, col_reg}<16'b1000110110110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110110110001) && ({row_reg, col_reg}<16'b1000110110110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110110110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000110110110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000110110110111) && ({row_reg, col_reg}<16'b1000110110111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000110110111001) && ({row_reg, col_reg}<16'b1000110110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110110111101) && ({row_reg, col_reg}<16'b1000110111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110111000000) && ({row_reg, col_reg}<16'b1000110111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000110111000011) && ({row_reg, col_reg}<16'b1000110111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110111000111) && ({row_reg, col_reg}<16'b1000110111001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000110111001010) && ({row_reg, col_reg}<16'b1000110111001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110111001100) && ({row_reg, col_reg}<16'b1000110111001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110111001111) && ({row_reg, col_reg}<16'b1000110111010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110111010001) && ({row_reg, col_reg}<16'b1000110111010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110111010101) && ({row_reg, col_reg}<16'b1000110111010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110111010111) && ({row_reg, col_reg}<16'b1000110111011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110111011100) && ({row_reg, col_reg}<16'b1000110111011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000110111011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000110111100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000110111100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000110111100010) && ({row_reg, col_reg}<16'b1000110111101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110111101010) && ({row_reg, col_reg}<16'b1000110111101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110111101101) && ({row_reg, col_reg}<16'b1000110111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110111110001) && ({row_reg, col_reg}<16'b1000110111110100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b1000110111110100) && ({row_reg, col_reg}<16'b1000111000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000111000000000) && ({row_reg, col_reg}<16'b1000111000000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111000000101) && ({row_reg, col_reg}<16'b1000111000000111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000111000000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1000111000001000)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==16'b1000111000001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000111000001010) && ({row_reg, col_reg}<16'b1000111000001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000111000001100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000111000001101) && ({row_reg, col_reg}<16'b1000111000001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111000001111) && ({row_reg, col_reg}<16'b1000111000010110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000111000010110) && ({row_reg, col_reg}<16'b1000111000011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111000011001) && ({row_reg, col_reg}<16'b1000111000011011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000111000011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111000011100) && ({row_reg, col_reg}<16'b1000111000011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111000011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000111000100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000111000100001) && ({row_reg, col_reg}<16'b1000111000100011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000111000100011) && ({row_reg, col_reg}<16'b1000111000101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000111000101001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000111000101010) && ({row_reg, col_reg}<16'b1000111000101110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111000101110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000111000101111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000111000110000) && ({row_reg, col_reg}<16'b1000111000110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111000110011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000111000110100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000111000110101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000111000110110) && ({row_reg, col_reg}<16'b1000111000111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111000111010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000111000111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000111000111100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000111000111101) && ({row_reg, col_reg}<16'b1000111001000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000111001000000) && ({row_reg, col_reg}<16'b1000111001000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000111001000010) && ({row_reg, col_reg}<16'b1000111001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111001000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111001000111) && ({row_reg, col_reg}<16'b1000111001001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111001001010) && ({row_reg, col_reg}<16'b1000111001001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000111001001100) && ({row_reg, col_reg}<16'b1000111001001110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1000111001001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000111001001111) && ({row_reg, col_reg}<16'b1000111001010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000111001010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000111001010110) && ({row_reg, col_reg}<16'b1000111001100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111001100110) && ({row_reg, col_reg}<16'b1000111001101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1000111001101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000111001101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000111001101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111001101101) && ({row_reg, col_reg}<16'b1000111001101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000111001101111) && ({row_reg, col_reg}<16'b1000111001110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111001110011) && ({row_reg, col_reg}<16'b1000111010000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111010000101) && ({row_reg, col_reg}<16'b1000111010001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111010001000) && ({row_reg, col_reg}<16'b1000111010001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111010001100) && ({row_reg, col_reg}<16'b1000111010001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111010001110) && ({row_reg, col_reg}<16'b1000111010010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000111010010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111010010001) && ({row_reg, col_reg}<16'b1000111010011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111010011101) && ({row_reg, col_reg}<16'b1000111010100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111010100000) && ({row_reg, col_reg}<16'b1000111010101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111010101010) && ({row_reg, col_reg}<16'b1000111010101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111010101100) && ({row_reg, col_reg}<16'b1000111010110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111010110001) && ({row_reg, col_reg}<16'b1000111010110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111010110011) && ({row_reg, col_reg}<16'b1000111010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000111010110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000111010110110) && ({row_reg, col_reg}<16'b1000111010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000111010111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000111010111001) && ({row_reg, col_reg}<16'b1000111010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000111010111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000111010111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111011000000) && ({row_reg, col_reg}<16'b1000111011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000111011000011) && ({row_reg, col_reg}<16'b1000111011000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111011000111) && ({row_reg, col_reg}<16'b1000111011001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000111011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111011001011) && ({row_reg, col_reg}<16'b1000111011010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111011010000) && ({row_reg, col_reg}<16'b1000111011010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111011010101) && ({row_reg, col_reg}<16'b1000111011011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111011011000) && ({row_reg, col_reg}<16'b1000111011011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111011011100) && ({row_reg, col_reg}<16'b1000111011011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111011011111) && ({row_reg, col_reg}<16'b1000111011100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000111011100011) && ({row_reg, col_reg}<16'b1000111011100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000111011100101) && ({row_reg, col_reg}<16'b1000111011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111011110001) && ({row_reg, col_reg}<16'b1000111011110100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b1000111011110100) && ({row_reg, col_reg}<16'b1000111100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000111100000000) && ({row_reg, col_reg}<16'b1000111100000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111100000101) && ({row_reg, col_reg}<16'b1000111100000111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000111100000111) && ({row_reg, col_reg}<16'b1000111100001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000111100001001) && ({row_reg, col_reg}<16'b1000111100001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000111100001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000111100001110) && ({row_reg, col_reg}<16'b1000111100010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111100010100) && ({row_reg, col_reg}<16'b1000111100010111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000111100010111) && ({row_reg, col_reg}<16'b1000111100011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000111100011011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000111100011100) && ({row_reg, col_reg}<16'b1000111100011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111100011110) && ({row_reg, col_reg}<16'b1000111100100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111100100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000111100100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111100100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000111100100011) && ({row_reg, col_reg}<16'b1000111100101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000111100101000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000111100101001) && ({row_reg, col_reg}<16'b1000111100101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111100101111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000111100110000) && ({row_reg, col_reg}<16'b1000111100110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111100110100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000111100110101) && ({row_reg, col_reg}<16'b1000111100111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000111100111010) && ({row_reg, col_reg}<16'b1000111101000000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000111101000000) && ({row_reg, col_reg}<16'b1000111101000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000111101000011) && ({row_reg, col_reg}<16'b1000111101000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000111101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000111101000111) && ({row_reg, col_reg}<16'b1000111101001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000111101001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000111101001010) && ({row_reg, col_reg}<16'b1000111101010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000111101010001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000111101010010) && ({row_reg, col_reg}<16'b1000111101010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000111101010100) && ({row_reg, col_reg}<16'b1000111101011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000111101011101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000111101011110) && ({row_reg, col_reg}<16'b1000111101100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111101100000) && ({row_reg, col_reg}<16'b1000111101100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000111101100100) && ({row_reg, col_reg}<16'b1000111101100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111101100110) && ({row_reg, col_reg}<16'b1000111101101000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b1000111101101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000111101101001) && ({row_reg, col_reg}<16'b1000111101101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000111101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000111101101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000111101101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000111101101110) && ({row_reg, col_reg}<16'b1000111101110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111101110001) && ({row_reg, col_reg}<16'b1000111110000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111110000110) && ({row_reg, col_reg}<16'b1000111110001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111110001001) && ({row_reg, col_reg}<16'b1000111110001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111110001011) && ({row_reg, col_reg}<16'b1000111110001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000111110001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111110001111) && ({row_reg, col_reg}<16'b1000111110010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111110010010) && ({row_reg, col_reg}<16'b1000111110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111110110000) && ({row_reg, col_reg}<16'b1000111110110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111110110010) && ({row_reg, col_reg}<16'b1000111110110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000111110110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111110110101) && ({row_reg, col_reg}<16'b1000111110111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000111110111011) && ({row_reg, col_reg}<16'b1000111111000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111111000000) && ({row_reg, col_reg}<16'b1000111111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000111111000011) && ({row_reg, col_reg}<16'b1000111111000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111111000110) && ({row_reg, col_reg}<16'b1000111111001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111111001100) && ({row_reg, col_reg}<16'b1000111111001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111111001111) && ({row_reg, col_reg}<16'b1000111111010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111111010110) && ({row_reg, col_reg}<16'b1000111111011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111111011000) && ({row_reg, col_reg}<16'b1000111111011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111111011101) && ({row_reg, col_reg}<16'b1000111111011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111111011111) && ({row_reg, col_reg}<16'b1000111111100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000111111100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000111111100110) && ({row_reg, col_reg}<16'b1000111111101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000111111101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000111111101001) && ({row_reg, col_reg}<16'b1000111111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111111110001) && ({row_reg, col_reg}<16'b1000111111110100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b1000111111110100) && ({row_reg, col_reg}<16'b1001000000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001000000000000) && ({row_reg, col_reg}<16'b1001000000000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001000000000010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b1001000000000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001000000000100) && ({row_reg, col_reg}<16'b1001000000000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001000000000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001000000000111) && ({row_reg, col_reg}<16'b1001000000001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000000001010) && ({row_reg, col_reg}<16'b1001000000001100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001000000001100) && ({row_reg, col_reg}<16'b1001000000010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000000010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001000000010011) && ({row_reg, col_reg}<16'b1001000000010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000000010101) && ({row_reg, col_reg}<16'b1001000000011001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001000000011001) && ({row_reg, col_reg}<16'b1001000000011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000000011100) && ({row_reg, col_reg}<16'b1001000000011110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001000000011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000000011111) && ({row_reg, col_reg}<16'b1001000000100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001000000100011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001000000100100) && ({row_reg, col_reg}<16'b1001000000100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001000000100111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1001000000101000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001000000101001) && ({row_reg, col_reg}<16'b1001000000101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001000000101111) && ({row_reg, col_reg}<16'b1001000000110001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001000000110001) && ({row_reg, col_reg}<16'b1001000001000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001000001000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000001000011) && ({row_reg, col_reg}<16'b1001000001001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001000001001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001000001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000001001100) && ({row_reg, col_reg}<16'b1001000001001110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001000001001110) && ({row_reg, col_reg}<16'b1001000001010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000001010001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001000001010010) && ({row_reg, col_reg}<16'b1001000001011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000001011101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1001000001011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000001011111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001000001100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000001100001) && ({row_reg, col_reg}<16'b1001000001101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001000001101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000001101001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001000001101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000001101011) && ({row_reg, col_reg}<16'b1001000001101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000001101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001000001101110) && ({row_reg, col_reg}<16'b1001000001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000001110000) && ({row_reg, col_reg}<16'b1001000001110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000001110010) && ({row_reg, col_reg}<16'b1001000001110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000001110100) && ({row_reg, col_reg}<16'b1001000001111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000001111111) && ({row_reg, col_reg}<16'b1001000010000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001000010000001) && ({row_reg, col_reg}<16'b1001000010000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000010000011) && ({row_reg, col_reg}<16'b1001000010000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000010000111) && ({row_reg, col_reg}<16'b1001000010010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000010010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000010010001) && ({row_reg, col_reg}<16'b1001000010010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000010010011) && ({row_reg, col_reg}<16'b1001000010010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000010010101) && ({row_reg, col_reg}<16'b1001000010011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000010011001) && ({row_reg, col_reg}<16'b1001000010101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000010101111) && ({row_reg, col_reg}<16'b1001000010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000010110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001000010110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000010111000) && ({row_reg, col_reg}<16'b1001000010111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001000010111011) && ({row_reg, col_reg}<16'b1001000011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000011000000) && ({row_reg, col_reg}<16'b1001000011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001000011000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000011000100) && ({row_reg, col_reg}<16'b1001000011011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000011011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000011011001) && ({row_reg, col_reg}<16'b1001000011011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000011011101) && ({row_reg, col_reg}<16'b1001000011011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000011011111) && ({row_reg, col_reg}<16'b1001000011101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001000011101001) && ({row_reg, col_reg}<16'b1001000011101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001000011101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000011101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000011101101) && ({row_reg, col_reg}<16'b1001000011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000011110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001000011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001000011110011)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b1001000011110100) && ({row_reg, col_reg}<16'b1001000100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001000100000000) && ({row_reg, col_reg}<16'b1001000100000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001000100000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001000100000101) && ({row_reg, col_reg}<16'b1001000100001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000100001010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001000100001011) && ({row_reg, col_reg}<16'b1001000100001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000100001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001000100001110) && ({row_reg, col_reg}<16'b1001000100010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000100010010) && ({row_reg, col_reg}<16'b1001000100010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001000100010100) && ({row_reg, col_reg}<16'b1001000100011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000100011000) && ({row_reg, col_reg}<16'b1001000100011011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001000100011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000100011100) && ({row_reg, col_reg}<16'b1001000100100000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001000100100000) && ({row_reg, col_reg}<16'b1001000100100010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001000100100010) && ({row_reg, col_reg}<16'b1001000100100100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001000100100100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1001000100100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001000100100110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001000100100111) && ({row_reg, col_reg}<16'b1001000100101010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001000100101010) && ({row_reg, col_reg}<16'b1001000100101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001000100101111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001000100110000) && ({row_reg, col_reg}<16'b1001000101000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001000101000000) && ({row_reg, col_reg}<16'b1001000101000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000101000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001000101000011) && ({row_reg, col_reg}<16'b1001000101000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000101000110) && ({row_reg, col_reg}<16'b1001000101001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001000101001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001000101001011) && ({row_reg, col_reg}<16'b1001000101001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000101001110) && ({row_reg, col_reg}<16'b1001000101010000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001000101010000) && ({row_reg, col_reg}<16'b1001000101010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000101010011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001000101010100) && ({row_reg, col_reg}<16'b1001000101010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000101010110) && ({row_reg, col_reg}<16'b1001000101011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001000101011000) && ({row_reg, col_reg}<16'b1001000101011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000101011010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001000101011011) && ({row_reg, col_reg}<16'b1001000101011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000101011111) && ({row_reg, col_reg}<16'b1001000101100001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001000101100001) && ({row_reg, col_reg}<16'b1001000101100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000101100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001000101100110)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==16'b1001000101100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001000101101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000101101001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001000101101010) && ({row_reg, col_reg}<16'b1001000101101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000101101100) && ({row_reg, col_reg}<16'b1001000101101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001000101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000101101111) && ({row_reg, col_reg}<16'b1001000101110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000101110001) && ({row_reg, col_reg}<16'b1001000101110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000101110100) && ({row_reg, col_reg}<16'b1001000101111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001000101111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000101111111) && ({row_reg, col_reg}<16'b1001000110000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001000110000010) && ({row_reg, col_reg}<16'b1001000110000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000110000100) && ({row_reg, col_reg}<16'b1001000110000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000110000111) && ({row_reg, col_reg}<16'b1001000110010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000110010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000110010001) && ({row_reg, col_reg}<16'b1001000110010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000110010011) && ({row_reg, col_reg}<16'b1001000110010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000110010101) && ({row_reg, col_reg}<16'b1001000110011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000110011010) && ({row_reg, col_reg}<16'b1001000110101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000110101110) && ({row_reg, col_reg}<16'b1001000110110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000110110101) && ({row_reg, col_reg}<16'b1001000110111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000110111010) && ({row_reg, col_reg}<16'b1001000110111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000110111100) && ({row_reg, col_reg}<16'b1001000111000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001000111000000) && ({row_reg, col_reg}<16'b1001000111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001000111000011) && ({row_reg, col_reg}<16'b1001000111001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000111001010) && ({row_reg, col_reg}<16'b1001000111001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000111001100) && ({row_reg, col_reg}<16'b1001000111010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000111010110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001000111010111) && ({row_reg, col_reg}<16'b1001000111011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000111011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000111011010) && ({row_reg, col_reg}<16'b1001000111011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000111011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001000111011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000111011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001000111100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000111100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001000111100010) && ({row_reg, col_reg}<16'b1001000111101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001000111101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001000111101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000111101101) && ({row_reg, col_reg}<16'b1001000111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000111110001) && ({row_reg, col_reg}<16'b1001000111110101)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b1001000111110101) && ({row_reg, col_reg}<16'b1001001000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001001000000000) && ({row_reg, col_reg}<16'b1001001000000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001001000000100) && ({row_reg, col_reg}<16'b1001001000001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001000001101) && ({row_reg, col_reg}<16'b1001001000001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001001000001111) && ({row_reg, col_reg}<16'b1001001000010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001000010001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001001000010010) && ({row_reg, col_reg}<16'b1001001000010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001000010101) && ({row_reg, col_reg}<16'b1001001000011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001001000011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001000011001) && ({row_reg, col_reg}<16'b1001001000100000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001001000100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001000100001) && ({row_reg, col_reg}<16'b1001001000100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001001000100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001000100100) && ({row_reg, col_reg}<16'b1001001000101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001001000101000) && ({row_reg, col_reg}<16'b1001001000101011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001001000101011) && ({row_reg, col_reg}<16'b1001001000110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001001000110110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001001000110111) && ({row_reg, col_reg}<16'b1001001000111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001001000111111) && ({row_reg, col_reg}<16'b1001001001000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001001000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001001001000010) && ({row_reg, col_reg}<16'b1001001001000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001001000101) && ({row_reg, col_reg}<16'b1001001001000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001001001000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001001001000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001001001001001) && ({row_reg, col_reg}<16'b1001001001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001001001011)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b1001001001001100) && ({row_reg, col_reg}<16'b1001001001001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001001001001110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001001001001111) && ({row_reg, col_reg}<16'b1001001001010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001001010001) && ({row_reg, col_reg}<16'b1001001001010100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001001001010100) && ({row_reg, col_reg}<16'b1001001001010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001001010110) && ({row_reg, col_reg}<16'b1001001001011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001001001011000) && ({row_reg, col_reg}<16'b1001001001011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001001011010) && ({row_reg, col_reg}<16'b1001001001011100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001001001011100) && ({row_reg, col_reg}<16'b1001001001100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001001100000) && ({row_reg, col_reg}<16'b1001001001100010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001001001100010) && ({row_reg, col_reg}<16'b1001001001100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001001100101) && ({row_reg, col_reg}<16'b1001001001101001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001001001101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001001001101010) && ({row_reg, col_reg}<16'b1001001001101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001001101100) && ({row_reg, col_reg}<16'b1001001001101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001001001101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001001101111) && ({row_reg, col_reg}<16'b1001001001110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001001110001) && ({row_reg, col_reg}<16'b1001001001110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001001110100) && ({row_reg, col_reg}<16'b1001001001111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001001111100) && ({row_reg, col_reg}<16'b1001001001111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001001111110) && ({row_reg, col_reg}<16'b1001001010000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001001010000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001010000100) && ({row_reg, col_reg}<16'b1001001010000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001010000110) && ({row_reg, col_reg}<16'b1001001010001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001010001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001010001110) && ({row_reg, col_reg}<16'b1001001010010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001010010011) && ({row_reg, col_reg}<16'b1001001010011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001010011000) && ({row_reg, col_reg}<16'b1001001010011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001010011010) && ({row_reg, col_reg}<16'b1001001010011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001010011100) && ({row_reg, col_reg}<16'b1001001010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001010011111) && ({row_reg, col_reg}<16'b1001001010100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001001010100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001010100010) && ({row_reg, col_reg}<16'b1001001010100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001010100101) && ({row_reg, col_reg}<16'b1001001010100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001010100111) && ({row_reg, col_reg}<16'b1001001010101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001010101101) && ({row_reg, col_reg}<16'b1001001010110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001010110011) && ({row_reg, col_reg}<16'b1001001010110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001001010110101) && ({row_reg, col_reg}<16'b1001001010111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001001010111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001010111100) && ({row_reg, col_reg}<16'b1001001011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001001011000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001001011000100) && ({row_reg, col_reg}<16'b1001001011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001011001010) && ({row_reg, col_reg}<16'b1001001011001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001001011001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001011001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001001011001111) && ({row_reg, col_reg}<16'b1001001011010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001011010110) && ({row_reg, col_reg}<16'b1001001011011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001001011011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001011011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001011011010) && ({row_reg, col_reg}<16'b1001001011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001011011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001001011100000) && ({row_reg, col_reg}<16'b1001001011100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001011100010) && ({row_reg, col_reg}<16'b1001001011100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001001011100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001011100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001001011100110) && ({row_reg, col_reg}<16'b1001001011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001001011101111) && ({row_reg, col_reg}<16'b1001001011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001011110001) && ({row_reg, col_reg}<16'b1001001011110101)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b1001001011110101) && ({row_reg, col_reg}<16'b1001001100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001001100000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001100000001)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}>=16'b1001001100000010) && ({row_reg, col_reg}<16'b1001001100000100)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==16'b1001001100000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001001100000101) && ({row_reg, col_reg}<16'b1001001100001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001100001000) && ({row_reg, col_reg}<16'b1001001100001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001001100001100) && ({row_reg, col_reg}<16'b1001001100010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001100010001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001001100010010) && ({row_reg, col_reg}<16'b1001001100010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001100010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001001100010101) && ({row_reg, col_reg}<16'b1001001100011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001100011001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001001100011010) && ({row_reg, col_reg}<16'b1001001100011101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001001100011101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001001100011110) && ({row_reg, col_reg}<16'b1001001100100000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001001100100000) && ({row_reg, col_reg}<16'b1001001100100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001100100011) && ({row_reg, col_reg}<16'b1001001100100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001001100100101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001001100100110) && ({row_reg, col_reg}<16'b1001001100101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001001100101001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1001001100101010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001001100101011) && ({row_reg, col_reg}<16'b1001001100101101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001001100101101) && ({row_reg, col_reg}<16'b1001001100111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001001100111101) && ({row_reg, col_reg}<16'b1001001100111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001100111111) && ({row_reg, col_reg}<16'b1001001101000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001001101000110) && ({row_reg, col_reg}<16'b1001001101001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001101001011)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b1001001101001100) && ({row_reg, col_reg}<16'b1001001101001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001001101001110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001001101001111) && ({row_reg, col_reg}<16'b1001001101010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001101010110) && ({row_reg, col_reg}<16'b1001001101011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001001101011000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001001101011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001101011010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001001101011011) && ({row_reg, col_reg}<16'b1001001101011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001101011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001001101011110) && ({row_reg, col_reg}<16'b1001001101100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001101100000) && ({row_reg, col_reg}<16'b1001001101100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001001101100011) && ({row_reg, col_reg}<16'b1001001101100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001101100110) && ({row_reg, col_reg}<16'b1001001101101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001001101101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001001101101001) && ({row_reg, col_reg}<16'b1001001101110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001101110100) && ({row_reg, col_reg}<16'b1001001101111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001101111100) && ({row_reg, col_reg}<16'b1001001101111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001101111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001001101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001110000000) && ({row_reg, col_reg}<16'b1001001110000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001001110000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001001110000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001110000110) && ({row_reg, col_reg}<16'b1001001110001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001001110001010) && ({row_reg, col_reg}<16'b1001001110001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001110001100) && ({row_reg, col_reg}<16'b1001001110001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001110001111) && ({row_reg, col_reg}<16'b1001001110010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001110010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001110010011) && ({row_reg, col_reg}<16'b1001001110010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001110010101) && ({row_reg, col_reg}<16'b1001001110011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001110011100) && ({row_reg, col_reg}<16'b1001001110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001110011111) && ({row_reg, col_reg}<16'b1001001110101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001110101101) && ({row_reg, col_reg}<16'b1001001110101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001110101111) && ({row_reg, col_reg}<16'b1001001110110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001001110110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001110110011) && ({row_reg, col_reg}<16'b1001001110110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001001110110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001001110110111) && ({row_reg, col_reg}<16'b1001001110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001110111101) && ({row_reg, col_reg}<16'b1001001111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001001111000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001001111000100) && ({row_reg, col_reg}<16'b1001001111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001111001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001001111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001111001010) && ({row_reg, col_reg}<16'b1001001111001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001111001101) && ({row_reg, col_reg}<16'b1001001111010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001111010110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001001111010111) && ({row_reg, col_reg}<16'b1001001111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001111011111) && ({row_reg, col_reg}<16'b1001001111100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001001111100001) && ({row_reg, col_reg}<16'b1001001111100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001111100110) && ({row_reg, col_reg}<16'b1001001111101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001001111101000) && ({row_reg, col_reg}<16'b1001001111101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001001111101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001001111110000)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b1001001111110001) && ({row_reg, col_reg}<16'b1001010000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001010000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010000000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001010000000010)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}>=16'b1001010000000011) && ({row_reg, col_reg}<16'b1001010000000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010000000101) && ({row_reg, col_reg}<16'b1001010000001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010000001000) && ({row_reg, col_reg}<16'b1001010000001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010000001010)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==16'b1001010000001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001010000001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010000001101) && ({row_reg, col_reg}<16'b1001010000010000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010000010000) && ({row_reg, col_reg}<16'b1001010000010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010000010010) && ({row_reg, col_reg}<16'b1001010000010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001010000010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010000010101) && ({row_reg, col_reg}<16'b1001010000011000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001010000011000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001010000011001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001010000011010) && ({row_reg, col_reg}<16'b1001010000011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010000011111) && ({row_reg, col_reg}<16'b1001010000100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010000100001) && ({row_reg, col_reg}<16'b1001010000100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010000100100) && ({row_reg, col_reg}<16'b1001010000100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001010000100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010000101000) && ({row_reg, col_reg}<16'b1001010000101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001010000101010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001010000101011) && ({row_reg, col_reg}<16'b1001010000101101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001010000101101) && ({row_reg, col_reg}<16'b1001010000111100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001010000111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001010000111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010000111110) && ({row_reg, col_reg}<16'b1001010001000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010001000011) && ({row_reg, col_reg}<16'b1001010001000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010001000111) && ({row_reg, col_reg}<16'b1001010001001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001010001001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001010001001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001010001001100) && ({row_reg, col_reg}<16'b1001010001001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010001001111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010001010000) && ({row_reg, col_reg}<16'b1001010001010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010001010110) && ({row_reg, col_reg}<16'b1001010001011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001010001011000) && ({row_reg, col_reg}<16'b1001010001011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010001011100) && ({row_reg, col_reg}<16'b1001010001011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001010001011110) && ({row_reg, col_reg}<16'b1001010001100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001010001100000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1001010001100001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010001100010) && ({row_reg, col_reg}<16'b1001010001100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010001100100) && ({row_reg, col_reg}<16'b1001010001100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001010001100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010001101000) && ({row_reg, col_reg}<16'b1001010001101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010001101100) && ({row_reg, col_reg}<16'b1001010001101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010001101110) && ({row_reg, col_reg}<16'b1001010001110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010001110001) && ({row_reg, col_reg}<16'b1001010001110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001010001110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010001110100) && ({row_reg, col_reg}<16'b1001010001111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010001111101) && ({row_reg, col_reg}<16'b1001010001111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010001111111) && ({row_reg, col_reg}<16'b1001010010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001010010000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010010000010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010010000011) && ({row_reg, col_reg}<16'b1001010010000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010010000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001010010001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010010001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010010001010) && ({row_reg, col_reg}<16'b1001010010010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010010010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010010010001) && ({row_reg, col_reg}<16'b1001010010010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010010010011) && ({row_reg, col_reg}<16'b1001010010010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010010010110) && ({row_reg, col_reg}<16'b1001010010011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010010011100) && ({row_reg, col_reg}<16'b1001010010011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010010011110) && ({row_reg, col_reg}<16'b1001010010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010010110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010010110011) && ({row_reg, col_reg}<16'b1001010010111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010010111000) && ({row_reg, col_reg}<16'b1001010010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010010111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010011000000) && ({row_reg, col_reg}<16'b1001010011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001010011000100) && ({row_reg, col_reg}<16'b1001010011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010011001010) && ({row_reg, col_reg}<16'b1001010011001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010011001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001010011001101) && ({row_reg, col_reg}<16'b1001010011011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010011011111) && ({row_reg, col_reg}<16'b1001010011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001010011100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001010011100010) && ({row_reg, col_reg}<16'b1001010011100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010011100111) && ({row_reg, col_reg}<16'b1001010011101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001010011101001) && ({row_reg, col_reg}<16'b1001010011101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001010011101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001010011101100) && ({row_reg, col_reg}<16'b1001010011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001010011101111) && ({row_reg, col_reg}<16'b1001010011110001)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b1001010011110001) && ({row_reg, col_reg}<16'b1001010100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001010100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010100000001) && ({row_reg, col_reg}<16'b1001010100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001010100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010100001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001010100001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001010100001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010100001101) && ({row_reg, col_reg}<16'b1001010100010000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001010100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010100010001) && ({row_reg, col_reg}<16'b1001010100010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010100010100) && ({row_reg, col_reg}<16'b1001010100010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010100010110) && ({row_reg, col_reg}<16'b1001010100011000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010100011000) && ({row_reg, col_reg}<16'b1001010100011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010100011010) && ({row_reg, col_reg}<16'b1001010100100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010100100000) && ({row_reg, col_reg}<16'b1001010100100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010100100010) && ({row_reg, col_reg}<16'b1001010100100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010100100101) && ({row_reg, col_reg}<16'b1001010100101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001010100101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010100101010) && ({row_reg, col_reg}<16'b1001010100110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001010100110000) && ({row_reg, col_reg}<16'b1001010100110101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001010100110101) && ({row_reg, col_reg}<16'b1001010100111100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001010100111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001010100111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010100111110) && ({row_reg, col_reg}<16'b1001010101000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010101000000) && ({row_reg, col_reg}<16'b1001010101000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010101000010) && ({row_reg, col_reg}<16'b1001010101000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010101000111) && ({row_reg, col_reg}<16'b1001010101001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001010101001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001010101001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001010101001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010101001101) && ({row_reg, col_reg}<16'b1001010101001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010101001111) && ({row_reg, col_reg}<16'b1001010101010001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010101010001) && ({row_reg, col_reg}<16'b1001010101010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001010101010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001010101011000) && ({row_reg, col_reg}<16'b1001010101011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010101011100) && ({row_reg, col_reg}<16'b1001010101011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001010101011110) && ({row_reg, col_reg}<16'b1001010101100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010101100010) && ({row_reg, col_reg}<16'b1001010101100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010101100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001010101100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001010101100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010101100111) && ({row_reg, col_reg}<16'b1001010101101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010101101100) && ({row_reg, col_reg}<16'b1001010101101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010101101110) && ({row_reg, col_reg}<16'b1001010101110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010101110011) && ({row_reg, col_reg}<16'b1001010101110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010101110101) && ({row_reg, col_reg}<16'b1001010101111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010101111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001010101111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010101111010) && ({row_reg, col_reg}<16'b1001010101111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001010101111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010101111110) && ({row_reg, col_reg}<16'b1001010110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001010110000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010110000011) && ({row_reg, col_reg}<16'b1001010110010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010110010010) && ({row_reg, col_reg}<16'b1001010110010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010110010110) && ({row_reg, col_reg}<16'b1001010110011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010110011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010110011111) && ({row_reg, col_reg}<16'b1001010110100001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010110100001) && ({row_reg, col_reg}<16'b1001010110100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010110100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001010110100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001010110100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010110100110) && ({row_reg, col_reg}<16'b1001010110101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010110101001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001010110101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010110101100) && ({row_reg, col_reg}<16'b1001010110101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010110101110) && ({row_reg, col_reg}<16'b1001010110110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010110110010) && ({row_reg, col_reg}<16'b1001010110110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010110110111) && ({row_reg, col_reg}<16'b1001010110111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010110111001) && ({row_reg, col_reg}<16'b1001010110111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010110111100) && ({row_reg, col_reg}<16'b1001010110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001010110111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010111000000)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=16'b1001010111000001) && ({row_reg, col_reg}<16'b1001010111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001010111000100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001010111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001010111000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001010111000111) && ({row_reg, col_reg}<16'b1001010111001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001010111001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001010111001101) && ({row_reg, col_reg}<16'b1001010111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010111011111) && ({row_reg, col_reg}<16'b1001010111100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001010111100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001010111100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001010111100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010111100100) && ({row_reg, col_reg}<16'b1001010111101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010111101011) && ({row_reg, col_reg}<16'b1001010111101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010111101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001010111101110) && ({row_reg, col_reg}<16'b1001010111110000)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b1001010111110000) && ({row_reg, col_reg}<16'b1001011000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001011000000000) && ({row_reg, col_reg}<16'b1001011000000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001011000000011) && ({row_reg, col_reg}<16'b1001011000010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011000010101) && ({row_reg, col_reg}<16'b1001011000010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001011000010111) && ({row_reg, col_reg}<16'b1001011000011001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001011000011001) && ({row_reg, col_reg}<16'b1001011000011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011000011101) && ({row_reg, col_reg}<16'b1001011000011111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011000011111) && ({row_reg, col_reg}<16'b1001011000100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011000100001) && ({row_reg, col_reg}<16'b1001011000100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011000100011) && ({row_reg, col_reg}<16'b1001011000100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011000100101) && ({row_reg, col_reg}<16'b1001011000101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001011000101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011000101011) && ({row_reg, col_reg}<16'b1001011000110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001011000110010) && ({row_reg, col_reg}<16'b1001011000110111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001011000110111) && ({row_reg, col_reg}<16'b1001011000111100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001011000111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001011000111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011000111110) && ({row_reg, col_reg}<16'b1001011001000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011001000000) && ({row_reg, col_reg}<16'b1001011001000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001011001000010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001011001000011) && ({row_reg, col_reg}<16'b1001011001001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001011001001000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001011001001001) && ({row_reg, col_reg}<16'b1001011001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011001001011) && ({row_reg, col_reg}<16'b1001011001001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001011001001111) && ({row_reg, col_reg}<16'b1001011001010001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001011001010001) && ({row_reg, col_reg}<16'b1001011001011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011001011100) && ({row_reg, col_reg}<16'b1001011001011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001011001011111) && ({row_reg, col_reg}<16'b1001011001100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011001100010) && ({row_reg, col_reg}<16'b1001011001100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001011001100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011001100110) && ({row_reg, col_reg}<16'b1001011001101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011001101100) && ({row_reg, col_reg}<16'b1001011001110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001011001110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011001110010) && ({row_reg, col_reg}<16'b1001011001111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011001111101) && ({row_reg, col_reg}<16'b1001011010000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011010000100) && ({row_reg, col_reg}<16'b1001011010010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011010010001) && ({row_reg, col_reg}<16'b1001011010010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011010010101) && ({row_reg, col_reg}<16'b1001011010011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001011010011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011010011111) && ({row_reg, col_reg}<16'b1001011010100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011010100110) && ({row_reg, col_reg}<16'b1001011010101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011010101001) && ({row_reg, col_reg}<16'b1001011010101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011010101110) && ({row_reg, col_reg}<16'b1001011010110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011010110001) && ({row_reg, col_reg}<16'b1001011010110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011010110111) && ({row_reg, col_reg}<16'b1001011010111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011010111010) && ({row_reg, col_reg}<16'b1001011010111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011010111101) && ({row_reg, col_reg}<16'b1001011010111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001011010111111) && ({row_reg, col_reg}<16'b1001011011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011011000001) && ({row_reg, col_reg}<16'b1001011011000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011011000011) && ({row_reg, col_reg}<16'b1001011011001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001011011001000) && ({row_reg, col_reg}<16'b1001011011011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011011011110) && ({row_reg, col_reg}<16'b1001011011100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001011011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001011011100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001011011100010) && ({row_reg, col_reg}<16'b1001011011101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011011101000) && ({row_reg, col_reg}<16'b1001011011101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001011011101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001011011110000)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=16'b1001011011110001) && ({row_reg, col_reg}<16'b1001011100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001011100000000) && ({row_reg, col_reg}<16'b1001011100000010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001011100000010) && ({row_reg, col_reg}<16'b1001011100010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011100010001) && ({row_reg, col_reg}<16'b1001011100010011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001011100010011) && ({row_reg, col_reg}<16'b1001011100010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011100010101) && ({row_reg, col_reg}<16'b1001011100010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001011100010111)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b1001011100011000) && ({row_reg, col_reg}<16'b1001011100011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001011100011010) && ({row_reg, col_reg}<16'b1001011100011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001011100011101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001011100011110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001011100011111) && ({row_reg, col_reg}<16'b1001011100100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011100100001) && ({row_reg, col_reg}<16'b1001011100100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011100100101) && ({row_reg, col_reg}<16'b1001011100101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011100101010) && ({row_reg, col_reg}<16'b1001011100101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011100101100) && ({row_reg, col_reg}<16'b1001011100101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011100101111) && ({row_reg, col_reg}<16'b1001011100110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001011100110010) && ({row_reg, col_reg}<16'b1001011100110100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001011100110100) && ({row_reg, col_reg}<16'b1001011100111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001011100111010) && ({row_reg, col_reg}<16'b1001011100111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011100111101) && ({row_reg, col_reg}<16'b1001011101000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011101000011) && ({row_reg, col_reg}<16'b1001011101001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011101001110) && ({row_reg, col_reg}<16'b1001011101010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001011101010000) && ({row_reg, col_reg}<16'b1001011101010010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001011101010010) && ({row_reg, col_reg}<16'b1001011101010100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001011101010100) && ({row_reg, col_reg}<16'b1001011101011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011101011100) && ({row_reg, col_reg}<16'b1001011101100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001011101100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011101100001) && ({row_reg, col_reg}<16'b1001011101100011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1001011101100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001011101100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001011101100101) && ({row_reg, col_reg}<16'b1001011101100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011101100111) && ({row_reg, col_reg}<16'b1001011101101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001011101101010) && ({row_reg, col_reg}<16'b1001011101101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001011101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001011101101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001011101101110) && ({row_reg, col_reg}<16'b1001011101110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001011101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011101110001) && ({row_reg, col_reg}<16'b1001011101111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011101111100) && ({row_reg, col_reg}<16'b1001011110000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011110000100) && ({row_reg, col_reg}<16'b1001011110001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001011110001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011110001100) && ({row_reg, col_reg}<16'b1001011110001111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001011110001111) && ({row_reg, col_reg}<16'b1001011110010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001011110010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001011110010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011110011000) && ({row_reg, col_reg}<16'b1001011110011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001011110011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011110011111) && ({row_reg, col_reg}<16'b1001011110100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011110100010) && ({row_reg, col_reg}<16'b1001011110101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011110101000) && ({row_reg, col_reg}<16'b1001011110101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011110101010) && ({row_reg, col_reg}<16'b1001011110101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011110101110) && ({row_reg, col_reg}<16'b1001011110110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011110110001) && ({row_reg, col_reg}<16'b1001011110111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011110111000) && ({row_reg, col_reg}<16'b1001011110111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011110111010) && ({row_reg, col_reg}<16'b1001011110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011110111101) && ({row_reg, col_reg}<16'b1001011110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001011110111111) && ({row_reg, col_reg}<16'b1001011111000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011111000001) && ({row_reg, col_reg}<16'b1001011111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011111000101) && ({row_reg, col_reg}<16'b1001011111001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001011111001101) && ({row_reg, col_reg}<16'b1001011111011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011111011100) && ({row_reg, col_reg}<16'b1001011111011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001011111011111) && ({row_reg, col_reg}<16'b1001011111100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001011111100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001011111100010) && ({row_reg, col_reg}<16'b1001011111101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011111101000) && ({row_reg, col_reg}<16'b1001011111110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001011111110000)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b1001011111110001) && ({row_reg, col_reg}<16'b1001100000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001100000000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001100000000001) && ({row_reg, col_reg}<16'b1001100000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100000001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001100000001010) && ({row_reg, col_reg}<16'b1001100000010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100000010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001100000010010) && ({row_reg, col_reg}<16'b1001100000010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100000010101) && ({row_reg, col_reg}<16'b1001100000010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001100000010111) && ({row_reg, col_reg}<16'b1001100000011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001100000011001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001100000011010) && ({row_reg, col_reg}<16'b1001100000100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100000100000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001100000100001) && ({row_reg, col_reg}<16'b1001100000100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001100000100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100000100100) && ({row_reg, col_reg}<16'b1001100000100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100000100110) && ({row_reg, col_reg}<16'b1001100000101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100000101010) && ({row_reg, col_reg}<16'b1001100000101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100000101110) && ({row_reg, col_reg}<16'b1001100000110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100000110000) && ({row_reg, col_reg}<16'b1001100000111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001100000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100000111001) && ({row_reg, col_reg}<16'b1001100000111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100000111011) && ({row_reg, col_reg}<16'b1001100000111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100000111101) && ({row_reg, col_reg}<16'b1001100001000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100001000011) && ({row_reg, col_reg}<16'b1001100001001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100001001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001100001001100) && ({row_reg, col_reg}<16'b1001100001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100001001111) && ({row_reg, col_reg}<16'b1001100001010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001100001010001) && ({row_reg, col_reg}<16'b1001100001010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100001010011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001100001010100) && ({row_reg, col_reg}<16'b1001100001011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100001011001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001100001011010) && ({row_reg, col_reg}<16'b1001100001011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100001011100) && ({row_reg, col_reg}<16'b1001100001100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001100001100000) && ({row_reg, col_reg}<16'b1001100001100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100001100010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1001100001100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100001100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001100001100101) && ({row_reg, col_reg}<16'b1001100001100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100001100111) && ({row_reg, col_reg}<16'b1001100001101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001100001101001) && ({row_reg, col_reg}<16'b1001100001101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100001101011) && ({row_reg, col_reg}<16'b1001100001101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100001101110) && ({row_reg, col_reg}<16'b1001100001110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100001110010) && ({row_reg, col_reg}<16'b1001100010000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100010000000) && ({row_reg, col_reg}<16'b1001100010000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100010000110) && ({row_reg, col_reg}<16'b1001100010010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100010010000) && ({row_reg, col_reg}<16'b1001100010010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100010010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100010010101) && ({row_reg, col_reg}<16'b1001100010011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100010011001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100010011010) && ({row_reg, col_reg}<16'b1001100010011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100010011111) && ({row_reg, col_reg}<16'b1001100010100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100010100001) && ({row_reg, col_reg}<16'b1001100010101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100010101000) && ({row_reg, col_reg}<16'b1001100010110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100010110100) && ({row_reg, col_reg}<16'b1001100010111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100010111000) && ({row_reg, col_reg}<16'b1001100010111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100010111010) && ({row_reg, col_reg}<16'b1001100010111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100010111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100010111110) && ({row_reg, col_reg}<16'b1001100011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001100011000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001100011000001) && ({row_reg, col_reg}<16'b1001100011000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100011000011) && ({row_reg, col_reg}<16'b1001100011000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100011000111) && ({row_reg, col_reg}<16'b1001100011001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001100011001001) && ({row_reg, col_reg}<16'b1001100011001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001100011001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001100011001101) && ({row_reg, col_reg}<16'b1001100011011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100011011110) && ({row_reg, col_reg}<16'b1001100011100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001100011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001100011100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001100011100010) && ({row_reg, col_reg}<16'b1001100011100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100011100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001100011100110) && ({row_reg, col_reg}<16'b1001100011101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100011101000) && ({row_reg, col_reg}<16'b1001100011101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100011101010) && ({row_reg, col_reg}<16'b1001100011101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100011101100) && ({row_reg, col_reg}<16'b1001100011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001100011110000)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b1001100011110001) && ({row_reg, col_reg}<16'b1001100100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001100100000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001100100000001) && ({row_reg, col_reg}<16'b1001100100001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100100001010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001100100001011) && ({row_reg, col_reg}<16'b1001100100010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100100010000) && ({row_reg, col_reg}<16'b1001100100010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001100100010010) && ({row_reg, col_reg}<16'b1001100100010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100100010111) && ({row_reg, col_reg}<16'b1001100100011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001100100011001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001100100011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100100011011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001100100011100) && ({row_reg, col_reg}<16'b1001100100100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100100100000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1001100100100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100100100010) && ({row_reg, col_reg}<16'b1001100100100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100100100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001100100100101) && ({row_reg, col_reg}<16'b1001100100110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001100100110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001100100110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100100110010) && ({row_reg, col_reg}<16'b1001100100110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001100100110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100100110111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001100100111000) && ({row_reg, col_reg}<16'b1001100100111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100100111011) && ({row_reg, col_reg}<16'b1001100100111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100100111101) && ({row_reg, col_reg}<16'b1001100101000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100101000010) && ({row_reg, col_reg}<16'b1001100101001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100101001010) && ({row_reg, col_reg}<16'b1001100101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001100101001100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001100101001101) && ({row_reg, col_reg}<16'b1001100101010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100101010001) && ({row_reg, col_reg}<16'b1001100101010011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001100101010011) && ({row_reg, col_reg}<16'b1001100101010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100101010111) && ({row_reg, col_reg}<16'b1001100101011001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001100101011001) && ({row_reg, col_reg}<16'b1001100101011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100101011110) && ({row_reg, col_reg}<16'b1001100101100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001100101100000) && ({row_reg, col_reg}<16'b1001100101100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100101100011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001100101100100) && ({row_reg, col_reg}<16'b1001100101101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100101101011) && ({row_reg, col_reg}<16'b1001100101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100101101110) && ({row_reg, col_reg}<16'b1001100101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100101111011) && ({row_reg, col_reg}<16'b1001100101111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100101111101) && ({row_reg, col_reg}<16'b1001100110000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100110000111) && ({row_reg, col_reg}<16'b1001100110010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100110010010) && ({row_reg, col_reg}<16'b1001100110011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100110011001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001100110011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100110011011) && ({row_reg, col_reg}<16'b1001100110011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100110011111) && ({row_reg, col_reg}<16'b1001100110100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100110100011) && ({row_reg, col_reg}<16'b1001100110100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100110100101) && ({row_reg, col_reg}<16'b1001100110110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100110110011) && ({row_reg, col_reg}<16'b1001100110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100110110101) && ({row_reg, col_reg}<16'b1001100110110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100110110111) && ({row_reg, col_reg}<16'b1001100110111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100110111010) && ({row_reg, col_reg}<16'b1001100110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100110111110) && ({row_reg, col_reg}<16'b1001100111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100111000000) && ({row_reg, col_reg}<16'b1001100111000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100111000101) && ({row_reg, col_reg}<16'b1001100111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100111001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001100111001001) && ({row_reg, col_reg}<16'b1001100111001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001100111001101) && ({row_reg, col_reg}<16'b1001100111010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001100111010000) && ({row_reg, col_reg}<16'b1001100111011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100111011110) && ({row_reg, col_reg}<16'b1001100111100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001100111100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001100111100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001100111100010) && ({row_reg, col_reg}<16'b1001100111101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100111101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100111101001) && ({row_reg, col_reg}<16'b1001100111101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100111101100) && ({row_reg, col_reg}<16'b1001100111110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001100111110000)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b1001100111110001) && ({row_reg, col_reg}<16'b1001101000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001101000000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101000000001) && ({row_reg, col_reg}<16'b1001101000010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101000010001) && ({row_reg, col_reg}<16'b1001101000010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001101000010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101000010110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001101000010111) && ({row_reg, col_reg}<16'b1001101000011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101000011001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001101000011010) && ({row_reg, col_reg}<16'b1001101000011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101000011101) && ({row_reg, col_reg}<16'b1001101000011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001101000011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101000100000) && ({row_reg, col_reg}<16'b1001101000100010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1001101000100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101000100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001101000100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001101000100101) && ({row_reg, col_reg}<16'b1001101000100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101000100111) && ({row_reg, col_reg}<16'b1001101000101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101000101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001101000101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101000110000) && ({row_reg, col_reg}<16'b1001101000110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101000110010) && ({row_reg, col_reg}<16'b1001101000110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101000110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001101000110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101000110110) && ({row_reg, col_reg}<16'b1001101000111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101000111011) && ({row_reg, col_reg}<16'b1001101000111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101000111101) && ({row_reg, col_reg}<16'b1001101000111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101000111111) && ({row_reg, col_reg}<16'b1001101001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101001001001) && ({row_reg, col_reg}<16'b1001101001001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001101001001111) && ({row_reg, col_reg}<16'b1001101001010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101001010010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001101001010011) && ({row_reg, col_reg}<16'b1001101001011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101001011011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001101001011100) && ({row_reg, col_reg}<16'b1001101001011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101001011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001101001011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101001100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001101001100001) && ({row_reg, col_reg}<16'b1001101001100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101001100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001101001100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001101001100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001101001100110) && ({row_reg, col_reg}<16'b1001101001101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101001101001) && ({row_reg, col_reg}<16'b1001101001101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101001101111) && ({row_reg, col_reg}<16'b1001101001110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101001110010) && ({row_reg, col_reg}<16'b1001101001110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001101001110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101001110110) && ({row_reg, col_reg}<16'b1001101001111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001101001111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101001111011) && ({row_reg, col_reg}<16'b1001101001111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101001111110) && ({row_reg, col_reg}<16'b1001101010000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101010000001) && ({row_reg, col_reg}<16'b1001101010000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101010000101) && ({row_reg, col_reg}<16'b1001101010001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101010001000) && ({row_reg, col_reg}<16'b1001101010010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101010010011) && ({row_reg, col_reg}<16'b1001101010010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101010010110) && ({row_reg, col_reg}<16'b1001101010011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101010011000) && ({row_reg, col_reg}<16'b1001101010011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101010011011) && ({row_reg, col_reg}<16'b1001101010011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101010011110) && ({row_reg, col_reg}<16'b1001101010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101010100011) && ({row_reg, col_reg}<16'b1001101010100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101010100101) && ({row_reg, col_reg}<16'b1001101010100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101010100111) && ({row_reg, col_reg}<16'b1001101010110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101010110011) && ({row_reg, col_reg}<16'b1001101010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101010110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101010110110) && ({row_reg, col_reg}<16'b1001101010111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101010111000) && ({row_reg, col_reg}<16'b1001101010111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101010111101) && ({row_reg, col_reg}<16'b1001101011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101011000000) && ({row_reg, col_reg}<16'b1001101011000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101011000011) && ({row_reg, col_reg}<16'b1001101011000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101011000111) && ({row_reg, col_reg}<16'b1001101011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101011001001) && ({row_reg, col_reg}<16'b1001101011001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101011001100) && ({row_reg, col_reg}<16'b1001101011001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001101011001110) && ({row_reg, col_reg}<16'b1001101011010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001101011010000) && ({row_reg, col_reg}<16'b1001101011011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101011011110) && ({row_reg, col_reg}<16'b1001101011100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001101011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001101011100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001101011100010) && ({row_reg, col_reg}<16'b1001101011101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001101011101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101011101001) && ({row_reg, col_reg}<16'b1001101011101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101011101100) && ({row_reg, col_reg}<16'b1001101011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101011110000)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b1001101011110001) && ({row_reg, col_reg}<16'b1001101100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001101100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001101100000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001101100000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101100000011) && ({row_reg, col_reg}<16'b1001101100000101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001101100000101) && ({row_reg, col_reg}<16'b1001101100010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101100010001) && ({row_reg, col_reg}<16'b1001101100010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001101100010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101100010110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001101100010111) && ({row_reg, col_reg}<16'b1001101100011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101100011001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001101100011010) && ({row_reg, col_reg}<16'b1001101100011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101100011111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001101100100000) && ({row_reg, col_reg}<16'b1001101100100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101100100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001101100100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001101100100101) && ({row_reg, col_reg}<16'b1001101100101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101100101000) && ({row_reg, col_reg}<16'b1001101100101010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001101100101010) && ({row_reg, col_reg}<16'b1001101100101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101100101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001101100101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101100110000) && ({row_reg, col_reg}<16'b1001101100111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001101100111010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001101100111011) && ({row_reg, col_reg}<16'b1001101100111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101100111101) && ({row_reg, col_reg}<16'b1001101101000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001101101000000) && ({row_reg, col_reg}<16'b1001101101000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101101000101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001101101000110) && ({row_reg, col_reg}<16'b1001101101001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101101001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101101001011) && ({row_reg, col_reg}<16'b1001101101010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001101101010001) && ({row_reg, col_reg}<16'b1001101101010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101101010011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001101101010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001101101010101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001101101010110) && ({row_reg, col_reg}<16'b1001101101011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101101011110) && ({row_reg, col_reg}<16'b1001101101100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001101101100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101101100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101101100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101101100100) && ({row_reg, col_reg}<16'b1001101101100110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001101101100110) && ({row_reg, col_reg}<16'b1001101101110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101101110001) && ({row_reg, col_reg}<16'b1001101101111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101101111010) && ({row_reg, col_reg}<16'b1001101101111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101101111100) && ({row_reg, col_reg}<16'b1001101110000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101110000000) && ({row_reg, col_reg}<16'b1001101110000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101110000100) && ({row_reg, col_reg}<16'b1001101110001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101110001000) && ({row_reg, col_reg}<16'b1001101110010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101110010100) && ({row_reg, col_reg}<16'b1001101110010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001101110010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101110010111) && ({row_reg, col_reg}<16'b1001101110100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101110100111) && ({row_reg, col_reg}<16'b1001101110110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101110110010) && ({row_reg, col_reg}<16'b1001101110110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001101110110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101110110101) && ({row_reg, col_reg}<16'b1001101110110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001101110110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101110111000) && ({row_reg, col_reg}<16'b1001101110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001101110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101110111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001101110111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101111000000) && ({row_reg, col_reg}<16'b1001101111000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101111000010) && ({row_reg, col_reg}<16'b1001101111000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001101111000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101111000101) && ({row_reg, col_reg}<16'b1001101111001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101111001000) && ({row_reg, col_reg}<16'b1001101111001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101111001100) && ({row_reg, col_reg}<16'b1001101111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101111001110) && ({row_reg, col_reg}<16'b1001101111010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001101111010011) && ({row_reg, col_reg}<16'b1001101111011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101111011110) && ({row_reg, col_reg}<16'b1001101111100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001101111100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001101111100001) && ({row_reg, col_reg}<16'b1001101111100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001101111100011) && ({row_reg, col_reg}<16'b1001101111100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101111100111) && ({row_reg, col_reg}<16'b1001101111101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101111101001) && ({row_reg, col_reg}<16'b1001101111101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101111101100) && ({row_reg, col_reg}<16'b1001101111110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101111110000)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b1001101111110001) && ({row_reg, col_reg}<16'b1001110000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001110000000000) && ({row_reg, col_reg}<16'b1001110000000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110000000011) && ({row_reg, col_reg}<16'b1001110000000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110000000101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001110000000110) && ({row_reg, col_reg}<16'b1001110000001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110000001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001110000001110) && ({row_reg, col_reg}<16'b1001110000010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110000010011) && ({row_reg, col_reg}<16'b1001110000010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001110000010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110000010110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001110000010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110000011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110000011001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001110000011010) && ({row_reg, col_reg}<16'b1001110000100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110000100010) && ({row_reg, col_reg}<16'b1001110000100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001110000100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110000100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001110000101000) && ({row_reg, col_reg}<16'b1001110000101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110000101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001110000101100) && ({row_reg, col_reg}<16'b1001110000101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110000101110) && ({row_reg, col_reg}<16'b1001110000110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001110000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110000110101) && ({row_reg, col_reg}<16'b1001110000110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110000110111) && ({row_reg, col_reg}<16'b1001110000111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110000111011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1001110000111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110000111101) && ({row_reg, col_reg}<16'b1001110001000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001110001000001) && ({row_reg, col_reg}<16'b1001110001000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110001000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001110001000100) && ({row_reg, col_reg}<16'b1001110001001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110001001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001110001001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001110001001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110001001101) && ({row_reg, col_reg}<16'b1001110001001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001110001001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110001010000) && ({row_reg, col_reg}<16'b1001110001010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001110001010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110001010011) && ({row_reg, col_reg}<16'b1001110001010110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110001010110) && ({row_reg, col_reg}<16'b1001110001011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110001011000) && ({row_reg, col_reg}<16'b1001110001011010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001110001011010) && ({row_reg, col_reg}<16'b1001110001011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110001011100) && ({row_reg, col_reg}<16'b1001110001100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001110001100000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001110001100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110001100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110001100011) && ({row_reg, col_reg}<16'b1001110001100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001110001100101) && ({row_reg, col_reg}<16'b1001110001101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110001101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110001101010) && ({row_reg, col_reg}<16'b1001110001101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110001101101) && ({row_reg, col_reg}<16'b1001110001110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110001110101) && ({row_reg, col_reg}<16'b1001110001110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110001110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110001111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110001111001) && ({row_reg, col_reg}<16'b1001110001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110001111011) && ({row_reg, col_reg}<16'b1001110001111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001110001111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110001111111) && ({row_reg, col_reg}<16'b1001110010000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110010000100) && ({row_reg, col_reg}<16'b1001110010001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110010001000) && ({row_reg, col_reg}<16'b1001110010010111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110010010111) && ({row_reg, col_reg}<16'b1001110010011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110010011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110010011010) && ({row_reg, col_reg}<16'b1001110010011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110010011101) && ({row_reg, col_reg}<16'b1001110010100000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110010100000) && ({row_reg, col_reg}<16'b1001110010100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110010100101) && ({row_reg, col_reg}<16'b1001110010101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110010101111) && ({row_reg, col_reg}<16'b1001110010110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110010110011) && ({row_reg, col_reg}<16'b1001110010110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110010110101) && ({row_reg, col_reg}<16'b1001110010111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110010111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110010111010) && ({row_reg, col_reg}<16'b1001110010111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110010111101) && ({row_reg, col_reg}<16'b1001110011000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110011000011) && ({row_reg, col_reg}<16'b1001110011000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110011000110) && ({row_reg, col_reg}<16'b1001110011001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110011001000) && ({row_reg, col_reg}<16'b1001110011001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001110011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110011001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001110011001100) && ({row_reg, col_reg}<16'b1001110011001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110011001110) && ({row_reg, col_reg}<16'b1001110011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110011010001) && ({row_reg, col_reg}<16'b1001110011010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001110011010101) && ({row_reg, col_reg}<16'b1001110011011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110011011110) && ({row_reg, col_reg}<16'b1001110011100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001110011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001110011100001) && ({row_reg, col_reg}<16'b1001110011100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001110011100011) && ({row_reg, col_reg}<16'b1001110011100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110011100111) && ({row_reg, col_reg}<16'b1001110011101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110011101001) && ({row_reg, col_reg}<16'b1001110011101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110011101100) && ({row_reg, col_reg}<16'b1001110011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110011110000)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b1001110011110001) && ({row_reg, col_reg}<16'b1001110100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001110100000000) && ({row_reg, col_reg}<16'b1001110100000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110100000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110100000101) && ({row_reg, col_reg}<16'b1001110100000111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001110100000111) && ({row_reg, col_reg}<16'b1001110100001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110100001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001110100001010) && ({row_reg, col_reg}<16'b1001110100001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110100001101) && ({row_reg, col_reg}<16'b1001110100001111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001110100001111) && ({row_reg, col_reg}<16'b1001110100010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110100010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001110100010101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001110100010110) && ({row_reg, col_reg}<16'b1001110100011000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110100011000) && ({row_reg, col_reg}<16'b1001110100011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001110100011010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001110100011011) && ({row_reg, col_reg}<16'b1001110100100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110100100100) && ({row_reg, col_reg}<16'b1001110100100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001110100100110) && ({row_reg, col_reg}<16'b1001110100101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110100101011) && ({row_reg, col_reg}<16'b1001110100101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001110100101101) && ({row_reg, col_reg}<16'b1001110100101111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001110100101111) && ({row_reg, col_reg}<16'b1001110100110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110100110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001110100110011) && ({row_reg, col_reg}<16'b1001110100110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110100110110) && ({row_reg, col_reg}<16'b1001110100111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110100111011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001110100111100) && ({row_reg, col_reg}<16'b1001110101000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110101000111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001110101001000) && ({row_reg, col_reg}<16'b1001110101001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110101001010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001110101001011) && ({row_reg, col_reg}<16'b1001110101001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110101001101) && ({row_reg, col_reg}<16'b1001110101001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001110101001111) && ({row_reg, col_reg}<16'b1001110101010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110101010001)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}>=16'b1001110101010010) && ({row_reg, col_reg}<16'b1001110101010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110101010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001110101010101) && ({row_reg, col_reg}<16'b1001110101011001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001110101011001) && ({row_reg, col_reg}<16'b1001110101011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110101011101) && ({row_reg, col_reg}<16'b1001110101011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001110101011111) && ({row_reg, col_reg}<16'b1001110101100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110101100001) && ({row_reg, col_reg}<16'b1001110101100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110101100011) && ({row_reg, col_reg}<16'b1001110101100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001110101100101) && ({row_reg, col_reg}<16'b1001110101101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110101101000) && ({row_reg, col_reg}<16'b1001110101110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001110101110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110101110100) && ({row_reg, col_reg}<16'b1001110101111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110101111000) && ({row_reg, col_reg}<16'b1001110101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110101111011) && ({row_reg, col_reg}<16'b1001110101111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110101111110) && ({row_reg, col_reg}<16'b1001110110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110110000000) && ({row_reg, col_reg}<16'b1001110110000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110110000010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001110110000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110110000100) && ({row_reg, col_reg}<16'b1001110110001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110110001011) && ({row_reg, col_reg}<16'b1001110110011000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001110110011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110110011001) && ({row_reg, col_reg}<16'b1001110110011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110110011011) && ({row_reg, col_reg}<16'b1001110110011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110110011101) && ({row_reg, col_reg}<16'b1001110110100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110110100001) && ({row_reg, col_reg}<16'b1001110110100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110110100011) && ({row_reg, col_reg}<16'b1001110110101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110110101000) && ({row_reg, col_reg}<16'b1001110110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110110101010) && ({row_reg, col_reg}<16'b1001110110101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001110110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110110101110) && ({row_reg, col_reg}<16'b1001110110110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110110110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110110110011) && ({row_reg, col_reg}<16'b1001110110110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110110110101) && ({row_reg, col_reg}<16'b1001110110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110110111101) && ({row_reg, col_reg}<16'b1001110110111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110110111111) && ({row_reg, col_reg}<16'b1001110111000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110111000010) && ({row_reg, col_reg}<16'b1001110111000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110111000100) && ({row_reg, col_reg}<16'b1001110111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110111000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001110111001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001110111001001) && ({row_reg, col_reg}<16'b1001110111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110111001011) && ({row_reg, col_reg}<16'b1001110111001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001110111001101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1001110111001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110111001111) && ({row_reg, col_reg}<16'b1001110111010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110111010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110111010011) && ({row_reg, col_reg}<16'b1001110111010110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001110111010110) && ({row_reg, col_reg}<16'b1001110111011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110111011110) && ({row_reg, col_reg}<16'b1001110111100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001110111100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001110111100001) && ({row_reg, col_reg}<16'b1001110111100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001110111100011) && ({row_reg, col_reg}<16'b1001110111101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110111101000) && ({row_reg, col_reg}<16'b1001110111101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110111101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110111101011) && ({row_reg, col_reg}<16'b1001110111101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110111101101) && ({row_reg, col_reg}<16'b1001110111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110111101111) && ({row_reg, col_reg}<16'b1001110111110001)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b1001110111110001) && ({row_reg, col_reg}<16'b1001111000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001111000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111000000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001111000000010) && ({row_reg, col_reg}<16'b1001111000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111000000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111000000111) && ({row_reg, col_reg}<16'b1001111000001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111000001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001111000001100) && ({row_reg, col_reg}<16'b1001111000001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111000001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001111000010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111000010001) && ({row_reg, col_reg}<16'b1001111000010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001111000010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111000010100) && ({row_reg, col_reg}<16'b1001111000010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001111000010110) && ({row_reg, col_reg}<16'b1001111000011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111000011000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001111000011001) && ({row_reg, col_reg}<16'b1001111000011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111000011100) && ({row_reg, col_reg}<16'b1001111000011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001111000011110) && ({row_reg, col_reg}<16'b1001111000100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111000100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001111000100001) && ({row_reg, col_reg}<16'b1001111000100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111000100100) && ({row_reg, col_reg}<16'b1001111000100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001111000100111) && ({row_reg, col_reg}<16'b1001111000101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111000101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001111000101101) && ({row_reg, col_reg}<16'b1001111000110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111000110000) && ({row_reg, col_reg}<16'b1001111000110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001111000110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111000110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001111000110100) && ({row_reg, col_reg}<16'b1001111000110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111000110110) && ({row_reg, col_reg}<16'b1001111000111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111000111000) && ({row_reg, col_reg}<16'b1001111000111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001111000111011) && ({row_reg, col_reg}<16'b1001111000111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111000111110) && ({row_reg, col_reg}<16'b1001111001000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001111001000000) && ({row_reg, col_reg}<16'b1001111001000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111001000011) && ({row_reg, col_reg}<16'b1001111001000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001111001000101) && ({row_reg, col_reg}<16'b1001111001001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111001001001) && ({row_reg, col_reg}<16'b1001111001001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001111001001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111001001101) && ({row_reg, col_reg}<16'b1001111001001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001111001001111) && ({row_reg, col_reg}<16'b1001111001010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111001010010) && ({row_reg, col_reg}<16'b1001111001010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001111001010101) && ({row_reg, col_reg}<16'b1001111001011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111001011001) && ({row_reg, col_reg}<16'b1001111001011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001111001011011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001111001011100) && ({row_reg, col_reg}<16'b1001111001011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111001011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111001100000) && ({row_reg, col_reg}<16'b1001111001100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111001100111) && ({row_reg, col_reg}<16'b1001111001110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001111001110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111001110100) && ({row_reg, col_reg}<16'b1001111001111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111001111001) && ({row_reg, col_reg}<16'b1001111010000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111010000011) && ({row_reg, col_reg}<16'b1001111010001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111010001011) && ({row_reg, col_reg}<16'b1001111010011000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111010011000) && ({row_reg, col_reg}<16'b1001111010011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111010011010) && ({row_reg, col_reg}<16'b1001111010011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111010011100) && ({row_reg, col_reg}<16'b1001111010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111010011111) && ({row_reg, col_reg}<16'b1001111010100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111010100111) && ({row_reg, col_reg}<16'b1001111010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111010101010) && ({row_reg, col_reg}<16'b1001111010101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001111010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111010101110) && ({row_reg, col_reg}<16'b1001111010110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001111010110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111010110010) && ({row_reg, col_reg}<16'b1001111010110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111010110101) && ({row_reg, col_reg}<16'b1001111010110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111010110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111010111000) && ({row_reg, col_reg}<16'b1001111010111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111010111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111010111110) && ({row_reg, col_reg}<16'b1001111011000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111011000010) && ({row_reg, col_reg}<16'b1001111011000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111011000100) && ({row_reg, col_reg}<16'b1001111011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111011001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111011001001) && ({row_reg, col_reg}<16'b1001111011001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111011001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111011001101) && ({row_reg, col_reg}<16'b1001111011001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111011001111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001111011010000) && ({row_reg, col_reg}<16'b1001111011010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111011010010) && ({row_reg, col_reg}<16'b1001111011011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111011011001) && ({row_reg, col_reg}<16'b1001111011011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001111011011100) && ({row_reg, col_reg}<16'b1001111011011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111011011110) && ({row_reg, col_reg}<16'b1001111011100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001111011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001111011100001) && ({row_reg, col_reg}<16'b1001111011100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001111011100011) && ({row_reg, col_reg}<16'b1001111011101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111011101000) && ({row_reg, col_reg}<16'b1001111011101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111011101101) && ({row_reg, col_reg}<16'b1001111011110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111011110000)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=16'b1001111011110001) && ({row_reg, col_reg}<16'b1001111100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001111100000000) && ({row_reg, col_reg}<16'b1001111100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111100000110) && ({row_reg, col_reg}<16'b1001111100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001111100001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001111100001001) && ({row_reg, col_reg}<16'b1001111100001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111100001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001111100001100) && ({row_reg, col_reg}<16'b1001111100001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111100001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001111100001111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b1001111100010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b1001111100010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001111100010010) && ({row_reg, col_reg}<16'b1001111100010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111100010100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b1001111100010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b1001111100010110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b1001111100010111) && ({row_reg, col_reg}<16'b1001111100011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111100011100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001111100011101) && ({row_reg, col_reg}<16'b1001111100011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001111100011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111100100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001111100100001) && ({row_reg, col_reg}<16'b1001111100100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111100100011) && ({row_reg, col_reg}<16'b1001111100100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001111100100101) && ({row_reg, col_reg}<16'b1001111100101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111100101000) && ({row_reg, col_reg}<16'b1001111100101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001111100101010) && ({row_reg, col_reg}<16'b1001111100110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111100110000) && ({row_reg, col_reg}<16'b1001111100110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001111100110011) && ({row_reg, col_reg}<16'b1001111100111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111100111000) && ({row_reg, col_reg}<16'b1001111100111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001111100111011) && ({row_reg, col_reg}<16'b1001111100111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111100111110) && ({row_reg, col_reg}<16'b1001111101000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001111101000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111101000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001111101000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111101000011) && ({row_reg, col_reg}<16'b1001111101000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001111101000110) && ({row_reg, col_reg}<16'b1001111101001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111101001000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001111101001001) && ({row_reg, col_reg}<16'b1001111101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001111101001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111101001101) && ({row_reg, col_reg}<16'b1001111101010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001111101010000) && ({row_reg, col_reg}<16'b1001111101010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111101010011) && ({row_reg, col_reg}<16'b1001111101010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001111101010110) && ({row_reg, col_reg}<16'b1001111101011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111101011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001111101011011) && ({row_reg, col_reg}<16'b1001111101011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111101011110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001111101011111) && ({row_reg, col_reg}<16'b1001111101100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111101100010) && ({row_reg, col_reg}<16'b1001111101100100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001111101100100) && ({row_reg, col_reg}<16'b1001111101100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111101100111) && ({row_reg, col_reg}<16'b1001111101110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111101110101) && ({row_reg, col_reg}<16'b1001111101111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111101111000) && ({row_reg, col_reg}<16'b1001111110000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111110000011) && ({row_reg, col_reg}<16'b1001111110000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111110000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111110000110) && ({row_reg, col_reg}<16'b1001111110001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111110001000) && ({row_reg, col_reg}<16'b1001111110001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111110001010) && ({row_reg, col_reg}<16'b1001111110001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111110001100) && ({row_reg, col_reg}<16'b1001111110001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111110001110) && ({row_reg, col_reg}<16'b1001111110011001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111110011001) && ({row_reg, col_reg}<16'b1001111110011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111110011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111110011111) && ({row_reg, col_reg}<16'b1001111110100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111110100001) && ({row_reg, col_reg}<16'b1001111110100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111110100111) && ({row_reg, col_reg}<16'b1001111110101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111110101110) && ({row_reg, col_reg}<16'b1001111110110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001111110110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111110110001) && ({row_reg, col_reg}<16'b1001111110110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111110110101) && ({row_reg, col_reg}<16'b1001111110111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111110111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001111110111011) && ({row_reg, col_reg}<16'b1001111111000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111111000010) && ({row_reg, col_reg}<16'b1001111111000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111111000100) && ({row_reg, col_reg}<16'b1001111111001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111111001100) && ({row_reg, col_reg}<16'b1001111111010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111111010011) && ({row_reg, col_reg}<16'b1001111111010101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001111111010101) && ({row_reg, col_reg}<16'b1001111111010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111111010111) && ({row_reg, col_reg}<16'b1001111111011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111111011001) && ({row_reg, col_reg}<16'b1001111111011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001111111011100) && ({row_reg, col_reg}<16'b1001111111011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111111011110) && ({row_reg, col_reg}<16'b1001111111100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001111111100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001111111100001) && ({row_reg, col_reg}<16'b1001111111100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001111111100011) && ({row_reg, col_reg}<16'b1001111111101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111111101000) && ({row_reg, col_reg}<16'b1001111111110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001111111110000)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=16'b1001111111110001) && ({row_reg, col_reg}<=16'b1001111111111111)) color_data = 12'b000000000000;
	end
endmodule