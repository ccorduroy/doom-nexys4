module bgl_rom
	(
		input wire clk,
		input wire [7:0] row,
		input wire [7:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [7:0] row_reg;
	reg [7:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin
		if(({row_reg, col_reg}==16'b0000000000000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000000000001) && ({row_reg, col_reg}<16'b0000000000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000000000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000000000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000000000000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0000000000001000) && ({row_reg, col_reg}<16'b0000000000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000000000001100) && ({row_reg, col_reg}<16'b0000000000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000000010000) && ({row_reg, col_reg}<16'b0000000000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000000010010) && ({row_reg, col_reg}<16'b0000000001100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000000001100010) && ({row_reg, col_reg}<16'b0000000001100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000001100111) && ({row_reg, col_reg}<16'b0000000001101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000000001101001) && ({row_reg, col_reg}<16'b0000000001101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000001101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000001101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000001101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000000001101111) && ({row_reg, col_reg}<16'b0000000001110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000001110001) && ({row_reg, col_reg}<16'b0000000001110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000000001110011) && ({row_reg, col_reg}<16'b0000000001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000001111101) && ({row_reg, col_reg}<16'b0000000010000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000010000010) && ({row_reg, col_reg}<16'b0000000010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000000010010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000010010101) && ({row_reg, col_reg}<16'b0000000010010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000010010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000010011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000010011001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000000010011010) && ({row_reg, col_reg}<16'b0000000010011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000010011101) && ({row_reg, col_reg}<16'b0000000010100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000010100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000010100001) && ({row_reg, col_reg}<16'b0000000010100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000000010100011) && ({row_reg, col_reg}<16'b0000000010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000000010100101) && ({row_reg, col_reg}<16'b0000000010100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000000010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000010101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000000010101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000010101010) && ({row_reg, col_reg}<16'b0000000010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000010110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000000010110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000000010110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000000010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000000010110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000010110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000000010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000010110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000000010111000) && ({row_reg, col_reg}<16'b0000000010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000000010111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000000010111011)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==16'b0000000010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000010111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000000010111110) && ({row_reg, col_reg}<16'b0000000011000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000011000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000000011000101) && ({row_reg, col_reg}<16'b0000000011000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000000011000111) && ({row_reg, col_reg}<16'b0000000011001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000000011001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000000011001100) && ({row_reg, col_reg}<16'b0000000011001110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000000011001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000011001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000000011010000) && ({row_reg, col_reg}<16'b0000000011010010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000000011010010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000000011010011) && ({row_reg, col_reg}<16'b0000000011010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000000011010101) && ({row_reg, col_reg}<16'b0000000011010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000011010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000000011011000) && ({row_reg, col_reg}<16'b0000000011011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000000011011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000011011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000000011011100) && ({row_reg, col_reg}<16'b0000000011011110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000000011011110) && ({row_reg, col_reg}<16'b0000000011100000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000011100000)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0000000011100001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000000011100010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000000011100011) && ({row_reg, col_reg}<16'b0000000011100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000011100101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000000011100110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000011100111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000000011101000)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0000000011101001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000000011101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000011101011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000000011101100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000011101101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000000011101110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000000011101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000011110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000011110001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000000011110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000011110011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000000011110100)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0000000011110101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000000011110110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000011110111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000000011111000) && ({row_reg, col_reg}<16'b0000000011111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000011111010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000000011111011) && ({row_reg, col_reg}<16'b0000000011111110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000000011111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0000000011111111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000000100000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000100000001) && ({row_reg, col_reg}<16'b0000000100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000100000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000000100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0000000100001000) && ({row_reg, col_reg}<16'b0000000100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000000100001100) && ({row_reg, col_reg}<16'b0000000100001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000100001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000000100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000100010000) && ({row_reg, col_reg}<16'b0000000100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000100010010) && ({row_reg, col_reg}<16'b0000000101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000000101100010) && ({row_reg, col_reg}<16'b0000000101100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000101100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000000101101000) && ({row_reg, col_reg}<16'b0000000101101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000101101011) && ({row_reg, col_reg}<16'b0000000101101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000101101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000101101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000000101101111) && ({row_reg, col_reg}<16'b0000000101110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000101110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000000101110010) && ({row_reg, col_reg}<16'b0000000101110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000101110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000000101110101) && ({row_reg, col_reg}<16'b0000000101111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000101111110) && ({row_reg, col_reg}<16'b0000000110000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000000110000010) && ({row_reg, col_reg}<16'b0000000110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000000110010100) && ({row_reg, col_reg}<16'b0000000110010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000110010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000110010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000110011000) && ({row_reg, col_reg}<16'b0000000110011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000000110011010) && ({row_reg, col_reg}<16'b0000000110011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000110011101) && ({row_reg, col_reg}<16'b0000000110100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000110100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000110100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000000110100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000000110100011) && ({row_reg, col_reg}<16'b0000000110100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000000110100111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0000000110101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000000110101001) && ({row_reg, col_reg}<16'b0000000110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000000110101101) && ({row_reg, col_reg}<16'b0000000110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000110110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000000110110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000000110110010) && ({row_reg, col_reg}<16'b0000000110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000000110110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000000110110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000000110110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000000110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000000110111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000000110111011) && ({row_reg, col_reg}<16'b0000000110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000000110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000000110111110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000110111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000000111000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000111000001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000000111000010) && ({row_reg, col_reg}<16'b0000000111000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000111000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000000111000101) && ({row_reg, col_reg}<16'b0000000111001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000000111001100) && ({row_reg, col_reg}<16'b0000000111001110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000000111001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000111001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000000111010000) && ({row_reg, col_reg}<16'b0000000111010010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000000111010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000000111010011) && ({row_reg, col_reg}<16'b0000000111010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000000111010101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000000111010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000111010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000000111011000) && ({row_reg, col_reg}<16'b0000000111011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000000111011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000000111011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000000111011100) && ({row_reg, col_reg}<16'b0000000111011110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000000111011110) && ({row_reg, col_reg}<16'b0000000111100000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000111100000)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0000000111100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000000111100010) && ({row_reg, col_reg}<16'b0000000111100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000111100111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000000111101000)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0000000111101001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000000111101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000111101011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000000111101100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000111101101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000000111101110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000000111101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000111110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000111110001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000000111110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000000111110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000000111110100) && ({row_reg, col_reg}<16'b0000000111110110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000000111110110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000000111110111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000000111111000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0000000111111001) && ({row_reg, col_reg}<16'b0000000111111011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000000111111011)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0000000111111100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0000000111111101)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0000000111111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0000000111111111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0000001000000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001000000001) && ({row_reg, col_reg}<16'b0000001000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001000000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000001000000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000001000001000) && ({row_reg, col_reg}<16'b0000001000001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000001000001011) && ({row_reg, col_reg}<16'b0000001000001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000001000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001000001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000001000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001000010000) && ({row_reg, col_reg}<16'b0000001000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001000010010) && ({row_reg, col_reg}<16'b0000001001100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000001001100010) && ({row_reg, col_reg}<16'b0000001001100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001001100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000001001101000) && ({row_reg, col_reg}<16'b0000001001101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001001101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000001001101100) && ({row_reg, col_reg}<16'b0000001001101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001001101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000001001101111) && ({row_reg, col_reg}<16'b0000001001110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001001110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000001001110010) && ({row_reg, col_reg}<16'b0000001001110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001001110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000001001110110) && ({row_reg, col_reg}<16'b0000001010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001010000010) && ({row_reg, col_reg}<16'b0000001010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000001010010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001010010101) && ({row_reg, col_reg}<16'b0000001010010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000001010010111) && ({row_reg, col_reg}<16'b0000001010011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001010011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000001010011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001010011101) && ({row_reg, col_reg}<16'b0000001010011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000001010011111) && ({row_reg, col_reg}<16'b0000001010100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001010100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000001010100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001010100011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000001010100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0000001010100101) && ({row_reg, col_reg}<16'b0000001010101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000001010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000001010101001) && ({row_reg, col_reg}<16'b0000001010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001010101101) && ({row_reg, col_reg}<16'b0000001010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000001010110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000001010110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000001010110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001010110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000001010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001010110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000001010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001010111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000001010111011) && ({row_reg, col_reg}<16'b0000001010111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000001010111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001010111110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000001010111111) && ({row_reg, col_reg}<16'b0000001011000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000001011000010) && ({row_reg, col_reg}<16'b0000001011001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000001011001100) && ({row_reg, col_reg}<16'b0000001011001110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000001011001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001011001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000001011010000) && ({row_reg, col_reg}<16'b0000001011010010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000001011010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001011010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001011010100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000001011010101) && ({row_reg, col_reg}<16'b0000001011010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000001011010111) && ({row_reg, col_reg}<16'b0000001011011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001011011001)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0000001011011010) && ({row_reg, col_reg}<16'b0000001011011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000001011011100) && ({row_reg, col_reg}<16'b0000001011011110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000001011011110) && ({row_reg, col_reg}<16'b0000001011100000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001011100000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000001011100001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000001011100010) && ({row_reg, col_reg}<16'b0000001011100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000001011100111) && ({row_reg, col_reg}<16'b0000001011101010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000001011101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001011101011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000001011101100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001011101101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000001011101110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000001011101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000001011110000) && ({row_reg, col_reg}<16'b0000001011110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000001011110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001011110011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000001011110100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000001011110101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0000001011110110) && ({row_reg, col_reg}<16'b0000001011111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001011111000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0000001011111001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000001011111010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000001011111011)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0000001011111100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0000001011111101)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0000001011111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0000001011111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000001100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000001100000001) && ({row_reg, col_reg}<16'b0000001100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001100000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000001100000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000001100001000) && ({row_reg, col_reg}<16'b0000001100001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000001100001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000001100001011) && ({row_reg, col_reg}<16'b0000001100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000001100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001100001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000001100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001100010000) && ({row_reg, col_reg}<16'b0000001100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001100010010) && ({row_reg, col_reg}<16'b0000001101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000001101100010) && ({row_reg, col_reg}<16'b0000001101100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001101100111) && ({row_reg, col_reg}<16'b0000001101101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000001101101001) && ({row_reg, col_reg}<16'b0000001101101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001101101101) && ({row_reg, col_reg}<16'b0000001101101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000001101101111) && ({row_reg, col_reg}<16'b0000001101110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001101110101) && ({row_reg, col_reg}<16'b0000001101110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000001101110111) && ({row_reg, col_reg}<16'b0000001110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000001110000010) && ({row_reg, col_reg}<16'b0000001110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000001110010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001110010101) && ({row_reg, col_reg}<16'b0000001110011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000001110011000) && ({row_reg, col_reg}<16'b0000001110011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001110011101) && ({row_reg, col_reg}<16'b0000001110011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000001110011111) && ({row_reg, col_reg}<16'b0000001110100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000001110100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000001110100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001110100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000001110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000001110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000001110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000001110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000001110101010) && ({row_reg, col_reg}<16'b0000001110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000001110110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000001110110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000001110110010) && ({row_reg, col_reg}<16'b0000001110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000001110110101) && ({row_reg, col_reg}<16'b0000001110111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000001110111000) && ({row_reg, col_reg}<16'b0000001110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000001110111011) && ({row_reg, col_reg}<16'b0000001110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000001110111110) && ({row_reg, col_reg}<16'b0000001111000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000001111000000) && ({row_reg, col_reg}<16'b0000001111000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000001111000010) && ({row_reg, col_reg}<16'b0000001111001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001111001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001111001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000001111010000) && ({row_reg, col_reg}<16'b0000001111010010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000001111010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000001111010011) && ({row_reg, col_reg}<16'b0000001111010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001111010110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000001111010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000001111011000) && ({row_reg, col_reg}<16'b0000001111011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000001111011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000001111011011) && ({row_reg, col_reg}<16'b0000001111011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000001111011110) && ({row_reg, col_reg}<16'b0000001111100010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000001111100010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001111100011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000001111100100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0000001111100101) && ({row_reg, col_reg}<16'b0000001111100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000001111100111) && ({row_reg, col_reg}<16'b0000001111101010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000001111101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001111101011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000001111101100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001111101101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000001111101110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000001111101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000001111110000) && ({row_reg, col_reg}<16'b0000001111110010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000001111110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001111110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001111110100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000001111110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000001111110110)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0000001111110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000001111111000)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0000001111111001)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0000001111111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000001111111011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000001111111100)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0000001111111101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000001111111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0000001111111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000010000000000) && ({row_reg, col_reg}<16'b0000010000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010000000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000010000000111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000010000001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000010000001010) && ({row_reg, col_reg}<16'b0000010000001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000010000001100) && ({row_reg, col_reg}<16'b0000010000001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010000001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010000001111) && ({row_reg, col_reg}<16'b0000010000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010000010010) && ({row_reg, col_reg}<16'b0000010001100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000010001100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010001100011) && ({row_reg, col_reg}<16'b0000010001101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010001101000) && ({row_reg, col_reg}<16'b0000010001101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000010001101010) && ({row_reg, col_reg}<16'b0000010001110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010001110101) && ({row_reg, col_reg}<16'b0000010001110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000010001110111) && ({row_reg, col_reg}<16'b0000010001111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010001111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000010001111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010001111011) && ({row_reg, col_reg}<16'b0000010001111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000010001111101) && ({row_reg, col_reg}<16'b0000010010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010010000010) && ({row_reg, col_reg}<16'b0000010010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000010010010100) && ({row_reg, col_reg}<16'b0000010010010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010010010110) && ({row_reg, col_reg}<16'b0000010010011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000010010011000) && ({row_reg, col_reg}<16'b0000010010100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010010100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000010010100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010010100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000010010100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000010010100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000010010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000010010100110) && ({row_reg, col_reg}<16'b0000010010101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000010010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000010010101001) && ({row_reg, col_reg}<16'b0000010010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000010010110000) && ({row_reg, col_reg}<16'b0000010010110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000010010110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000010010110011) && ({row_reg, col_reg}<16'b0000010010110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000010010110110) && ({row_reg, col_reg}<16'b0000010010111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000010010111000) && ({row_reg, col_reg}<16'b0000010010111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010010111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010010111100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0000010010111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000010010111110) && ({row_reg, col_reg}<16'b0000010011001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010011001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000010011001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010011001111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000010011010000) && ({row_reg, col_reg}<16'b0000010011010010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000010011010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000010011010011) && ({row_reg, col_reg}<16'b0000010011010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010011010101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000010011010110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010011010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000010011011000) && ({row_reg, col_reg}<16'b0000010011011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010011011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000010011011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010011011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000010011011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010011011110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000010011011111) && ({row_reg, col_reg}<16'b0000010011100010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010011100010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0000010011100011) && ({row_reg, col_reg}<16'b0000010011100101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0000010011100101) && ({row_reg, col_reg}<16'b0000010011100111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0000010011100111) && ({row_reg, col_reg}<16'b0000010011101010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000010011101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010011101011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000010011101100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000010011101101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000010011101110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000010011101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000010011110000) && ({row_reg, col_reg}<16'b0000010011110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000010011110010) && ({row_reg, col_reg}<16'b0000010011110100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010011110100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000010011110101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000010011110110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000010011110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010011111000) && ({row_reg, col_reg}<16'b0000010011111010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000010011111010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000010011111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010011111100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000010011111101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010011111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0000010011111111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0000010100000000) && ({row_reg, col_reg}<16'b0000010100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000010100000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000010100000111) && ({row_reg, col_reg}<16'b0000010100001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000010100001010) && ({row_reg, col_reg}<16'b0000010100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010100010010) && ({row_reg, col_reg}<16'b0000010101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000010101100010) && ({row_reg, col_reg}<16'b0000010101110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010101110100) && ({row_reg, col_reg}<16'b0000010101110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000010101110110) && ({row_reg, col_reg}<16'b0000010101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010101111000) && ({row_reg, col_reg}<16'b0000010101111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010101111010) && ({row_reg, col_reg}<16'b0000010101111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010101111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000010101111101) && ({row_reg, col_reg}<16'b0000010110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000010110000010) && ({row_reg, col_reg}<16'b0000010110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000010110010100) && ({row_reg, col_reg}<16'b0000010110010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010110010111) && ({row_reg, col_reg}<16'b0000010110011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000010110011011) && ({row_reg, col_reg}<16'b0000010110100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000010110100001) && ({row_reg, col_reg}<16'b0000010110100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000010110100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000010110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000010110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000010110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000010110101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000010110101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000010110101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000010110101101) && ({row_reg, col_reg}<16'b0000010110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000010110110000) && ({row_reg, col_reg}<16'b0000010110110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000010110110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000010110110011) && ({row_reg, col_reg}<16'b0000010110110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000010110110110) && ({row_reg, col_reg}<16'b0000010110111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000010110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000010110111001) && ({row_reg, col_reg}<16'b0000010110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010110111011) && ({row_reg, col_reg}<16'b0000010110111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000010110111111) && ({row_reg, col_reg}<16'b0000010111000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010111000111) && ({row_reg, col_reg}<16'b0000010111001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000010111001001) && ({row_reg, col_reg}<16'b0000010111001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010111001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000010111001110) && ({row_reg, col_reg}<16'b0000010111010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010111010000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010111010001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000010111010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000010111010011) && ({row_reg, col_reg}<16'b0000010111010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010111010110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000010111010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000010111011000) && ({row_reg, col_reg}<16'b0000010111011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000010111011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000010111011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010111011100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000010111011101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000010111011110) && ({row_reg, col_reg}<16'b0000010111100000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000010111100000) && ({row_reg, col_reg}<16'b0000010111101010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000010111101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010111101011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000010111101100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010111101101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000010111101110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000010111101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000010111110000) && ({row_reg, col_reg}<16'b0000010111110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010111110010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000010111110011) && ({row_reg, col_reg}<16'b0000010111110101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000010111110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000010111110110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000010111110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000010111111000) && ({row_reg, col_reg}<16'b0000010111111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000010111111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000010111111100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000010111111101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000010111111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0000010111111111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0000011000000000) && ({row_reg, col_reg}<16'b0000011000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011000000110) && ({row_reg, col_reg}<16'b0000011000001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000011000001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000011000001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011000001010) && ({row_reg, col_reg}<16'b0000011000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011000010010) && ({row_reg, col_reg}<16'b0000011001100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000011001100010) && ({row_reg, col_reg}<16'b0000011001110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011001110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000011001110101) && ({row_reg, col_reg}<16'b0000011001111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011001111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011001111010) && ({row_reg, col_reg}<16'b0000011010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011010000001) && ({row_reg, col_reg}<16'b0000011010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000011010010100) && ({row_reg, col_reg}<16'b0000011010010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011010010110) && ({row_reg, col_reg}<16'b0000011010011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011010011010) && ({row_reg, col_reg}<16'b0000011010100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011010100001) && ({row_reg, col_reg}<16'b0000011010100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000011010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000011010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000011010100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000011010101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000011010101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011010101010) && ({row_reg, col_reg}<16'b0000011010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011010110000) && ({row_reg, col_reg}<16'b0000011010110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000011010110011) && ({row_reg, col_reg}<16'b0000011010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000011010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000011010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000011010110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000011010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000011010111001) && ({row_reg, col_reg}<16'b0000011010111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000011010111011) && ({row_reg, col_reg}<16'b0000011010111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000011010111111) && ({row_reg, col_reg}<16'b0000011011000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000011011000111) && ({row_reg, col_reg}<16'b0000011011001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000011011001001) && ({row_reg, col_reg}<16'b0000011011001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000011011001101) && ({row_reg, col_reg}<16'b0000011011010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000011011010000) && ({row_reg, col_reg}<16'b0000011011010011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000011011010011) && ({row_reg, col_reg}<16'b0000011011011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000011011011000) && ({row_reg, col_reg}<16'b0000011011011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011011011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000011011011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000011011011100) && ({row_reg, col_reg}<16'b0000011011011111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000011011011111) && ({row_reg, col_reg}<16'b0000011011100010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011011100010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0000011011100011) && ({row_reg, col_reg}<16'b0000011011100110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0000011011100110) && ({row_reg, col_reg}<16'b0000011011101011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011011101011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000011011101100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011011101101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000011011101110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000011011101111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000011011110000) && ({row_reg, col_reg}<16'b0000011011110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011011110010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000011011110011) && ({row_reg, col_reg}<16'b0000011011110101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000011011110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011011110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011011110111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000011011111000) && ({row_reg, col_reg}<16'b0000011011111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011011111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011011111100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000011011111101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011011111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0000011011111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011100000001) && ({row_reg, col_reg}<16'b0000011100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011100000110) && ({row_reg, col_reg}<16'b0000011100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000011100001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000011100001001) && ({row_reg, col_reg}<16'b0000011100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011100001101) && ({row_reg, col_reg}<16'b0000011100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011100010010) && ({row_reg, col_reg}<16'b0000011101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000011101100010) && ({row_reg, col_reg}<16'b0000011101101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011101101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000011101101001) && ({row_reg, col_reg}<16'b0000011101101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011101101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000011101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011101101111) && ({row_reg, col_reg}<16'b0000011101110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011101110100) && ({row_reg, col_reg}<16'b0000011101110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011101110110) && ({row_reg, col_reg}<16'b0000011101111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011101111000) && ({row_reg, col_reg}<16'b0000011110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000011110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000011110000001) && ({row_reg, col_reg}<16'b0000011110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000011110010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011110010101) && ({row_reg, col_reg}<16'b0000011110011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000011110011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000011110011001) && ({row_reg, col_reg}<16'b0000011110011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000011110011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011110011101) && ({row_reg, col_reg}<16'b0000011110011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011110011111) && ({row_reg, col_reg}<16'b0000011110100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011110100011) && ({row_reg, col_reg}<16'b0000011110100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000011110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000011110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000011110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000011110101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000011110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000011110101010) && ({row_reg, col_reg}<16'b0000011110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000011110110000) && ({row_reg, col_reg}<16'b0000011110110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000011110110011) && ({row_reg, col_reg}<16'b0000011110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000011110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000011110110110) && ({row_reg, col_reg}<16'b0000011110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000011110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000011110111001) && ({row_reg, col_reg}<16'b0000011110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000011110111011) && ({row_reg, col_reg}<16'b0000011110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000011110111110) && ({row_reg, col_reg}<16'b0000011111000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000011111000110) && ({row_reg, col_reg}<16'b0000011111001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000011111001001) && ({row_reg, col_reg}<16'b0000011111001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011111001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000011111001101) && ({row_reg, col_reg}<16'b0000011111010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011111010000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000011111010001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011111010010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000011111010011) && ({row_reg, col_reg}<16'b0000011111010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011111010111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000011111011000) && ({row_reg, col_reg}<16'b0000011111011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000011111011010) && ({row_reg, col_reg}<16'b0000011111011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011111011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000011111011101) && ({row_reg, col_reg}<16'b0000011111011111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000011111011111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000011111100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011111100001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000011111100010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011111100011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000011111100100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0000011111100101) && ({row_reg, col_reg}<16'b0000011111101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011111101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000011111110000) && ({row_reg, col_reg}<16'b0000011111110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000011111110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011111110011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0000011111110100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000011111110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000011111110110) && ({row_reg, col_reg}<16'b0000011111111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000011111111010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000011111111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000011111111100) && ({row_reg, col_reg}<16'b0000011111111110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000011111111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0000011111111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000100000000000) && ({row_reg, col_reg}<16'b0000100000000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100000000010) && ({row_reg, col_reg}<16'b0000100000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100000000110) && ({row_reg, col_reg}<16'b0000100000001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000100000001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100000001011) && ({row_reg, col_reg}<16'b0000100000001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100000001101) && ({row_reg, col_reg}<16'b0000100000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100000010010) && ({row_reg, col_reg}<16'b0000100001100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000100001100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100001100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100001100100) && ({row_reg, col_reg}<16'b0000100001101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100001101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000100001101110) && ({row_reg, col_reg}<16'b0000100001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100001110000) && ({row_reg, col_reg}<16'b0000100001110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100001110100) && ({row_reg, col_reg}<16'b0000100001110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100001110110) && ({row_reg, col_reg}<16'b0000100001111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100001111000) && ({row_reg, col_reg}<16'b0000100010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100010000001) && ({row_reg, col_reg}<16'b0000100010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000100010010100) && ({row_reg, col_reg}<16'b0000100010010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100010010110) && ({row_reg, col_reg}<16'b0000100010011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100010011000) && ({row_reg, col_reg}<16'b0000100010011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000100010011101) && ({row_reg, col_reg}<16'b0000100010011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000100010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100010100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100010100001) && ({row_reg, col_reg}<16'b0000100010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100010100011) && ({row_reg, col_reg}<16'b0000100010100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000100010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000100010100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000100010101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000100010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100010101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000100010101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000100010101101) && ({row_reg, col_reg}<16'b0000100010101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000100010101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100010110000) && ({row_reg, col_reg}<16'b0000100010110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000100010110011) && ({row_reg, col_reg}<16'b0000100010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000100010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000100010110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000100010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100010111001) && ({row_reg, col_reg}<16'b0000100010111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000100010111011) && ({row_reg, col_reg}<16'b0000100010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100010111110) && ({row_reg, col_reg}<16'b0000100011000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100011000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100011000011) && ({row_reg, col_reg}<16'b0000100011000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000100011000110) && ({row_reg, col_reg}<16'b0000100011001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100011001001) && ({row_reg, col_reg}<16'b0000100011001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100011001100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000100011001101) && ({row_reg, col_reg}<16'b0000100011010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100011010000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100011010001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000100011010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100011010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000100011010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000100011010101) && ({row_reg, col_reg}<16'b0000100011010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000100011010111) && ({row_reg, col_reg}<16'b0000100011011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100011011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100011011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000100011011011) && ({row_reg, col_reg}<16'b0000100011100000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000100011100000) && ({row_reg, col_reg}<16'b0000100011100010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000100011100010) && ({row_reg, col_reg}<16'b0000100011100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100011100111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0000100011101000) && ({row_reg, col_reg}<16'b0000100011101011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000100011101011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0000100011101100) && ({row_reg, col_reg}<16'b0000100011101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100011101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100011110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100011110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000100011110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100011110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100011110100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000100011110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100011110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100011110111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000100011111000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100011111001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000100011111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100011111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100011111100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100011111101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000100011111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0000100011111111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0000100100000000) && ({row_reg, col_reg}<16'b0000100100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100100000010) && ({row_reg, col_reg}<16'b0000100100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100100000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000100100000111) && ({row_reg, col_reg}<16'b0000100100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000100100001001) && ({row_reg, col_reg}<16'b0000100100001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000100100001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000100100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100100001101) && ({row_reg, col_reg}<16'b0000100100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100100010010) && ({row_reg, col_reg}<16'b0000100101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000100101100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100101100011) && ({row_reg, col_reg}<16'b0000100101101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100101101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000100101101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100101101011) && ({row_reg, col_reg}<16'b0000100101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100101110000) && ({row_reg, col_reg}<16'b0000100101110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000100101110010) && ({row_reg, col_reg}<16'b0000100101111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100101111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000100101111101) && ({row_reg, col_reg}<16'b0000100110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100110000001) && ({row_reg, col_reg}<16'b0000100110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000100110010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100110010101) && ({row_reg, col_reg}<16'b0000100110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000100110010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100110011000) && ({row_reg, col_reg}<16'b0000100110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000100110011101) && ({row_reg, col_reg}<16'b0000100110011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000100110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100110100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000100110100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100110100010) && ({row_reg, col_reg}<16'b0000100110100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000100110100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000100110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000100110100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000100110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000100110101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000100110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000100110101011) && ({row_reg, col_reg}<16'b0000100110101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000100110101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000100110101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000100110101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0000100110110000) && ({row_reg, col_reg}<16'b0000100110110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100110110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000100110110011) && ({row_reg, col_reg}<16'b0000100110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000100110110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000100110110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000100110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100110111001) && ({row_reg, col_reg}<16'b0000100110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000100110111011) && ({row_reg, col_reg}<16'b0000100110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100110111101) && ({row_reg, col_reg}<16'b0000100110111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100110111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000100111000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100111000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100111000010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0000100111000011) && ({row_reg, col_reg}<16'b0000100111001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000100111001010) && ({row_reg, col_reg}<16'b0000100111001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100111001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000100111001110) && ({row_reg, col_reg}<16'b0000100111010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100111010000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100111010001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000100111010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100111010011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000100111010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000100111010101) && ({row_reg, col_reg}<16'b0000100111010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100111010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000100111011000) && ({row_reg, col_reg}<16'b0000100111011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100111011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000100111011011) && ({row_reg, col_reg}<16'b0000100111100000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000100111100000) && ({row_reg, col_reg}<16'b0000100111100010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000100111100010) && ({row_reg, col_reg}<16'b0000100111100110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100111100110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0000100111100111) && ({row_reg, col_reg}<16'b0000100111101100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000100111101100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000100111101101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000100111101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100111101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100111110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000100111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000100111110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000100111110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100111110100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000100111110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100111110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100111110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100111111000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100111111001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000100111111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000100111111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000100111111100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000100111111101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000100111111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0000100111111111)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0000101000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000101000000001) && ({row_reg, col_reg}<16'b0000101000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101000000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000101000000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000101000001000) && ({row_reg, col_reg}<16'b0000101000001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000101000001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000101000001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000101000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000101000001101) && ({row_reg, col_reg}<16'b0000101000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101000010010) && ({row_reg, col_reg}<16'b0000101001100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000101001100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101001100011) && ({row_reg, col_reg}<16'b0000101001101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101001101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000101001101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101001101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000101001101011) && ({row_reg, col_reg}<16'b0000101001101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101001101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000101001110000) && ({row_reg, col_reg}<16'b0000101001110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101001110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000101001110101) && ({row_reg, col_reg}<16'b0000101001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101001111111) && ({row_reg, col_reg}<16'b0000101010000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000101010000001) && ({row_reg, col_reg}<16'b0000101010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000101010010100) && ({row_reg, col_reg}<16'b0000101010010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000101010010111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101010011000) && ({row_reg, col_reg}<16'b0000101010011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000101010011101) && ({row_reg, col_reg}<16'b0000101010011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000101010011111) && ({row_reg, col_reg}<16'b0000101010100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101010100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000101010100010) && ({row_reg, col_reg}<16'b0000101010100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000101010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101010100110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000101010100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000101010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000101010101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000101010101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000101010101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101010101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000101010101101) && ({row_reg, col_reg}<16'b0000101010101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000101010101111) && ({row_reg, col_reg}<16'b0000101010110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0000101010110001) && ({row_reg, col_reg}<16'b0000101010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000101010110110) && ({row_reg, col_reg}<16'b0000101010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000101010111000) && ({row_reg, col_reg}<16'b0000101010111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101010111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101010111100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0000101010111101) && ({row_reg, col_reg}<16'b0000101010111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101010111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000101011000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101011000001) && ({row_reg, col_reg}<16'b0000101011000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000101011000101) && ({row_reg, col_reg}<16'b0000101011000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000101011000111) && ({row_reg, col_reg}<16'b0000101011001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000101011001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000101011001010) && ({row_reg, col_reg}<16'b0000101011001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101011001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000101011001110) && ({row_reg, col_reg}<16'b0000101011010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000101011010000) && ({row_reg, col_reg}<16'b0000101011010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101011010010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000101011010011) && ({row_reg, col_reg}<16'b0000101011010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101011010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000101011011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101011011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101011011010) && ({row_reg, col_reg}<16'b0000101011011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000101011011100) && ({row_reg, col_reg}<16'b0000101011100000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000101011100000) && ({row_reg, col_reg}<16'b0000101011100010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000101011100010) && ({row_reg, col_reg}<16'b0000101011100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101011100101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0000101011100110) && ({row_reg, col_reg}<16'b0000101011101100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000101011101100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000101011101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101011101110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101011101111) && ({row_reg, col_reg}<16'b0000101011110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000101011110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101011110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101011110011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000101011110100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000101011110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101011110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101011110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101011111000) && ({row_reg, col_reg}<16'b0000101011111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101011111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101011111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000101011111100) && ({row_reg, col_reg}<16'b0000101011111110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101011111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0000101011111111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000101100000000) && ({row_reg, col_reg}<16'b0000101100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101100000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000101100000111) && ({row_reg, col_reg}<16'b0000101100001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000101100001010) && ({row_reg, col_reg}<16'b0000101100001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000101100001100) && ({row_reg, col_reg}<16'b0000101100010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101100010011) && ({row_reg, col_reg}<16'b0000101100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000101100110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101100110101) && ({row_reg, col_reg}<16'b0000101100110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000101100110111) && ({row_reg, col_reg}<16'b0000101100111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000101100111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000101100111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101101000000) && ({row_reg, col_reg}<16'b0000101101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000101101011011) && ({row_reg, col_reg}<16'b0000101101011110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101101011110) && ({row_reg, col_reg}<16'b0000101101100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000101101100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000101101100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101101100010) && ({row_reg, col_reg}<16'b0000101101100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000101101100100) && ({row_reg, col_reg}<16'b0000101101100111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101101100111) && ({row_reg, col_reg}<16'b0000101101101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101101101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000101101101010) && ({row_reg, col_reg}<16'b0000101101101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000101101110000) && ({row_reg, col_reg}<16'b0000101101110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101101110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000101101110101) && ({row_reg, col_reg}<16'b0000101101111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101101111110) && ({row_reg, col_reg}<16'b0000101110000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000101110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101110000001) && ({row_reg, col_reg}<16'b0000101110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000101110010100) && ({row_reg, col_reg}<16'b0000101110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000101110010111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000101110011000) && ({row_reg, col_reg}<16'b0000101110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000101110011101) && ({row_reg, col_reg}<16'b0000101110011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000101110011111) && ({row_reg, col_reg}<16'b0000101110100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101110100010) && ({row_reg, col_reg}<16'b0000101110100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000101110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101110100110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000101110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000101110101000) && ({row_reg, col_reg}<16'b0000101110101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000101110101011) && ({row_reg, col_reg}<16'b0000101110101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000101110101101) && ({row_reg, col_reg}<16'b0000101110101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000101110101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0000101110110000) && ({row_reg, col_reg}<16'b0000101110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101110110011)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}==16'b0000101110110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000101110110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000101110110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000101110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000101110111001) && ({row_reg, col_reg}<16'b0000101110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101110111011) && ({row_reg, col_reg}<16'b0000101110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000101110111110) && ({row_reg, col_reg}<16'b0000101111000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101111000010) && ({row_reg, col_reg}<16'b0000101111000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101111000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000101111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000101111000110) && ({row_reg, col_reg}<16'b0000101111001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000101111001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000101111001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000101111001010) && ({row_reg, col_reg}<16'b0000101111001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101111001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000101111001110) && ({row_reg, col_reg}<16'b0000101111010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000101111010000) && ({row_reg, col_reg}<16'b0000101111010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101111010010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000101111010011) && ({row_reg, col_reg}<16'b0000101111010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101111010110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000101111010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000101111011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000101111011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101111011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000101111011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101111011100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000101111011101) && ({row_reg, col_reg}<16'b0000101111100000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101111100000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000101111100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101111100010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0000101111100011) && ({row_reg, col_reg}<16'b0000101111100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101111100101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0000101111100110) && ({row_reg, col_reg}<16'b0000101111101100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000101111101100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000101111101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101111101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000101111101111) && ({row_reg, col_reg}<16'b0000101111110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000101111110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101111110011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000101111110100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000101111110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101111110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101111110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000101111111000) && ({row_reg, col_reg}<16'b0000101111111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000101111111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000101111111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000101111111100) && ({row_reg, col_reg}<16'b0000101111111110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000101111111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0000101111111111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000110000000000) && ({row_reg, col_reg}<16'b0000110000000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110000000111) && ({row_reg, col_reg}<16'b0000110000001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000110000001010) && ({row_reg, col_reg}<16'b0000110000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110000010001) && ({row_reg, col_reg}<16'b0000110000010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000110000010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110000010100) && ({row_reg, col_reg}<16'b0000110000010110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110000010110) && ({row_reg, col_reg}<16'b0000110000011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110000011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110000011001) && ({row_reg, col_reg}<16'b0000110000011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000110000011011) && ({row_reg, col_reg}<16'b0000110000100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110000100000) && ({row_reg, col_reg}<16'b0000110000110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000110000110000) && ({row_reg, col_reg}<16'b0000110000110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110000110011) && ({row_reg, col_reg}<16'b0000110001000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110001000000) && ({row_reg, col_reg}<16'b0000110001000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110001000010) && ({row_reg, col_reg}<16'b0000110001010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000110001010111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000110001011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110001011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110001011010) && ({row_reg, col_reg}<16'b0000110001011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110001011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110001100000) && ({row_reg, col_reg}<16'b0000110001100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110001100010) && ({row_reg, col_reg}<16'b0000110001100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000110001100101) && ({row_reg, col_reg}<16'b0000110001101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110001101000) && ({row_reg, col_reg}<16'b0000110001101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000110001101010) && ({row_reg, col_reg}<16'b0000110001101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110001101100) && ({row_reg, col_reg}<16'b0000110001101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000110001101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110001101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000110001110000) && ({row_reg, col_reg}<16'b0000110001110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110001110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000110001110101) && ({row_reg, col_reg}<16'b0000110001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110001111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000110010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110010000001) && ({row_reg, col_reg}<16'b0000110010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000110010010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110010010101) && ({row_reg, col_reg}<16'b0000110010010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000110010010111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110010011000) && ({row_reg, col_reg}<16'b0000110010011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000110010011101) && ({row_reg, col_reg}<16'b0000110010011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000110010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110010100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110010100001) && ({row_reg, col_reg}<16'b0000110010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110010100011) && ({row_reg, col_reg}<16'b0000110010100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000110010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110010100110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000110010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110010101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000110010101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000110010101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000110010101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110010101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000110010101110) && ({row_reg, col_reg}<16'b0000110010110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110010110000) && ({row_reg, col_reg}<16'b0000110010110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000110010110010) && ({row_reg, col_reg}<16'b0000110010110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110010110110) && ({row_reg, col_reg}<16'b0000110010111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000110010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110010111001) && ({row_reg, col_reg}<16'b0000110010111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000110010111011) && ({row_reg, col_reg}<16'b0000110010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110010111110) && ({row_reg, col_reg}<16'b0000110011000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110011000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110011000011) && ({row_reg, col_reg}<16'b0000110011000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000110011000110) && ({row_reg, col_reg}<16'b0000110011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110011001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000110011001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110011001011) && ({row_reg, col_reg}<16'b0000110011001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000110011001110) && ({row_reg, col_reg}<16'b0000110011010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110011010000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000110011010001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000110011010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110011010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000110011010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110011010101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000110011010110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000110011010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110011011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110011011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110011011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000110011011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110011011100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000110011011101) && ({row_reg, col_reg}<16'b0000110011100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110011100001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000110011100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000110011100011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000110011100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110011100101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0000110011100110) && ({row_reg, col_reg}<16'b0000110011101100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000110011101100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000110011101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110011101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110011101111) && ({row_reg, col_reg}<16'b0000110011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110011110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110011110011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000110011110100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000110011110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110011110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110011110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000110011111000) && ({row_reg, col_reg}<16'b0000110011111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110011111010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000110011111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000110011111100) && ({row_reg, col_reg}<16'b0000110011111110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110011111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0000110011111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000110100000000) && ({row_reg, col_reg}<16'b0000110100000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110100000111) && ({row_reg, col_reg}<16'b0000110100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000110100001001) && ({row_reg, col_reg}<16'b0000110100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000110100001011) && ({row_reg, col_reg}<16'b0000110100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110100001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000110100001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110100001111) && ({row_reg, col_reg}<16'b0000110100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000110100010010) && ({row_reg, col_reg}<16'b0000110100011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110100011001) && ({row_reg, col_reg}<16'b0000110100011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110100011011) && ({row_reg, col_reg}<16'b0000110100011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110100011111) && ({row_reg, col_reg}<16'b0000110100101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110100101111) && ({row_reg, col_reg}<16'b0000110101000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110101000001) && ({row_reg, col_reg}<16'b0000110101010111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110101010111) && ({row_reg, col_reg}<16'b0000110101100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110101100001) && ({row_reg, col_reg}<16'b0000110101100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000110101100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110101100100) && ({row_reg, col_reg}<16'b0000110101100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000110101100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110101101000) && ({row_reg, col_reg}<16'b0000110101101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000110101101010) && ({row_reg, col_reg}<16'b0000110101101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110101101100) && ({row_reg, col_reg}<16'b0000110101101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000110101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000110101110000) && ({row_reg, col_reg}<16'b0000110101110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110101110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000110101110101) && ({row_reg, col_reg}<16'b0000110110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000110110000001) && ({row_reg, col_reg}<16'b0000110110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000110110010100) && ({row_reg, col_reg}<16'b0000110110011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110110011000) && ({row_reg, col_reg}<16'b0000110110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000110110011101) && ({row_reg, col_reg}<16'b0000110110011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000110110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110110100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000110110100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000110110100010) && ({row_reg, col_reg}<16'b0000110110100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000110110100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000110110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000110110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000110110101001) && ({row_reg, col_reg}<16'b0000110110110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000110110110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000110110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110110110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110110110110) && ({row_reg, col_reg}<16'b0000110110111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000110110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110110111001) && ({row_reg, col_reg}<16'b0000110110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110110111011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0000110110111100) && ({row_reg, col_reg}<16'b0000110110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110110111110) && ({row_reg, col_reg}<16'b0000110111000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110111000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110111000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000110111000100) && ({row_reg, col_reg}<16'b0000110111000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000110111000110) && ({row_reg, col_reg}<16'b0000110111001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000110111001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110111001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000110111001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000110111001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000110111001100) && ({row_reg, col_reg}<16'b0000110111001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110111001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110111001111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000110111010000) && ({row_reg, col_reg}<16'b0000110111010010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000110111010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110111010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000110111010100) && ({row_reg, col_reg}<16'b0000110111010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110111010110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000110111010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000110111011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000110111011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000110111011010) && ({row_reg, col_reg}<16'b0000110111011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0000110111011100) && ({row_reg, col_reg}<16'b0000110111011110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110111011110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0000110111011111) && ({row_reg, col_reg}<16'b0000110111101010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000110111101010)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0000110111101011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110111101100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000110111101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110111101110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000110111101111) && ({row_reg, col_reg}<16'b0000110111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000110111110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000110111110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000110111110011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000110111110100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0000110111110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110111110110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0000110111110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000110111111000) && ({row_reg, col_reg}<16'b0000110111111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000110111111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000110111111100) && ({row_reg, col_reg}<16'b0000110111111110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000110111111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0000110111111111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000111000000000) && ({row_reg, col_reg}<16'b0000111000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111000000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000111000000110) && ({row_reg, col_reg}<16'b0000111000001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111000001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000111000001001) && ({row_reg, col_reg}<16'b0000111000001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111000001110) && ({row_reg, col_reg}<16'b0000111000010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111000010011) && ({row_reg, col_reg}<16'b0000111000011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111000011000) && ({row_reg, col_reg}<16'b0000111000100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111000100011) && ({row_reg, col_reg}<16'b0000111000101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111000101001) && ({row_reg, col_reg}<16'b0000111000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111000110000) && ({row_reg, col_reg}<16'b0000111001000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111001000000) && ({row_reg, col_reg}<16'b0000111001011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111001011110) && ({row_reg, col_reg}<16'b0000111001100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111001100000) && ({row_reg, col_reg}<16'b0000111001100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111001100010) && ({row_reg, col_reg}<16'b0000111001100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111001100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000111001100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111001100110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000111001100111) && ({row_reg, col_reg}<16'b0000111001101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000111001101001) && ({row_reg, col_reg}<16'b0000111001110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111001110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000111001110101) && ({row_reg, col_reg}<16'b0000111010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111010000001) && ({row_reg, col_reg}<16'b0000111010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000111010010100) && ({row_reg, col_reg}<16'b0000111010010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111010010110) && ({row_reg, col_reg}<16'b0000111010011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000111010011000) && ({row_reg, col_reg}<16'b0000111010011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000111010011101) && ({row_reg, col_reg}<16'b0000111010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111010011111) && ({row_reg, col_reg}<16'b0000111010100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111010100001) && ({row_reg, col_reg}<16'b0000111010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111010100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111010100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000111010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000111010100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0000111010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000111010101001) && ({row_reg, col_reg}<16'b0000111010101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111010101110) && ({row_reg, col_reg}<16'b0000111010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111010110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000111010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111010110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000111010110101) && ({row_reg, col_reg}<16'b0000111010110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111010110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000111010111000) && ({row_reg, col_reg}<16'b0000111010111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000111010111011) && ({row_reg, col_reg}<16'b0000111010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000111010111110) && ({row_reg, col_reg}<16'b0000111011000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111011000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111011000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000111011000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111011000101) && ({row_reg, col_reg}<16'b0000111011001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000111011001001) && ({row_reg, col_reg}<16'b0000111011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111011001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000111011001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111011001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111011001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111011001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000111011010000) && ({row_reg, col_reg}<16'b0000111011010010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000111011010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000111011010011) && ({row_reg, col_reg}<16'b0000111011010101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000111011010101) && ({row_reg, col_reg}<16'b0000111011010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111011010111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0000111011011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111011011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000111011011010) && ({row_reg, col_reg}<16'b0000111011011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111011011100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000111011011101) && ({row_reg, col_reg}<16'b0000111011011111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000111011011111) && ({row_reg, col_reg}<16'b0000111011100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0000111011100010) && ({row_reg, col_reg}<16'b0000111011101000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0000111011101000) && ({row_reg, col_reg}<16'b0000111011101010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000111011101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111011101011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111011101100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111011101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111011101110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111011101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000111011110000) && ({row_reg, col_reg}<16'b0000111011110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111011110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111011110011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000111011110100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0000111011110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111011110110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0000111011110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111011111000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0000111011111001) && ({row_reg, col_reg}<16'b0000111011111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111011111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000111011111100) && ({row_reg, col_reg}<16'b0000111011111110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111011111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0000111011111111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0000111100000000) && ({row_reg, col_reg}<16'b0000111100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111100000110) && ({row_reg, col_reg}<16'b0000111100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111100001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0000111100001001) && ({row_reg, col_reg}<16'b0000111100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000111100001100) && ({row_reg, col_reg}<16'b0000111100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111100001111) && ({row_reg, col_reg}<16'b0000111100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111100010011) && ({row_reg, col_reg}<16'b0000111100010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000111100010110) && ({row_reg, col_reg}<16'b0000111100011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111100011010) && ({row_reg, col_reg}<16'b0000111100100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111100100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111100100010) && ({row_reg, col_reg}<16'b0000111100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000111100101010) && ({row_reg, col_reg}<16'b0000111100101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000111100101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111100101111) && ({row_reg, col_reg}<16'b0000111100110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111100110001) && ({row_reg, col_reg}<16'b0000111100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000111100110011) && ({row_reg, col_reg}<16'b0000111100110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111100110110) && ({row_reg, col_reg}<16'b0000111100111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000111100111000) && ({row_reg, col_reg}<16'b0000111100111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111100111010) && ({row_reg, col_reg}<16'b0000111100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000111100111101) && ({row_reg, col_reg}<16'b0000111101000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111101000001) && ({row_reg, col_reg}<16'b0000111101001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111101001010) && ({row_reg, col_reg}<16'b0000111101001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111101001110) && ({row_reg, col_reg}<16'b0000111101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000111101010000) && ({row_reg, col_reg}<16'b0000111101010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111101010101) && ({row_reg, col_reg}<16'b0000111101010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111101010111) && ({row_reg, col_reg}<16'b0000111101011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111101011001) && ({row_reg, col_reg}<16'b0000111101011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111101011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111101011110) && ({row_reg, col_reg}<16'b0000111101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000111101100001) && ({row_reg, col_reg}<16'b0000111101100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111101100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000111101100101) && ({row_reg, col_reg}<16'b0000111101100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000111101100111) && ({row_reg, col_reg}<16'b0000111101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000111101101011) && ({row_reg, col_reg}<16'b0000111101110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111101110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000111101110101) && ({row_reg, col_reg}<16'b0000111110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111110000001) && ({row_reg, col_reg}<16'b0000111110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0000111110010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111110010101) && ({row_reg, col_reg}<16'b0000111110011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0000111110011000) && ({row_reg, col_reg}<16'b0000111110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000111110011101) && ({row_reg, col_reg}<16'b0000111110100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111110100000) && ({row_reg, col_reg}<16'b0000111110100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0000111110100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111110100011) && ({row_reg, col_reg}<16'b0000111110100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0000111110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111110101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0000111110101001) && ({row_reg, col_reg}<16'b0000111110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0000111110101101) && ({row_reg, col_reg}<16'b0000111110110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111110110001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0000111110110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000111110110011) && ({row_reg, col_reg}<16'b0000111110110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000111110110110) && ({row_reg, col_reg}<16'b0000111110111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111110111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111110111001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000111110111010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0000111110111011) && ({row_reg, col_reg}<16'b0000111110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0000111110111101) && ({row_reg, col_reg}<16'b0000111111000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111111000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111111000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111111000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111111000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0000111111000110) && ({row_reg, col_reg}<16'b0000111111001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0000111111001010) && ({row_reg, col_reg}<16'b0000111111001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0000111111001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111111001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111111001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111111001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000111111010000) && ({row_reg, col_reg}<16'b0000111111010010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0000111111010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000111111010011) && ({row_reg, col_reg}<16'b0000111111010101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0000111111010101) && ({row_reg, col_reg}<16'b0000111111010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111111010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111111011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111111011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000111111011010) && ({row_reg, col_reg}<16'b0000111111011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111111011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000111111011101) && ({row_reg, col_reg}<16'b0000111111011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111111011111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000111111100000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000111111100001) && ({row_reg, col_reg}<16'b0000111111100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111111100011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000111111100100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000111111100101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0000111111100110) && ({row_reg, col_reg}<16'b0000111111101011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0000111111101011) && ({row_reg, col_reg}<16'b0000111111101101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0000111111101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111111101110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000111111101111) && ({row_reg, col_reg}<16'b0000111111110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0000111111110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0000111111110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111111110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0000111111110100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111111110101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0000111111110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0000111111110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0000111111111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0000111111111001) && ({row_reg, col_reg}<16'b0000111111111011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0000111111111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0000111111111100) && ({row_reg, col_reg}<16'b0000111111111110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0000111111111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0000111111111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001000000000000) && ({row_reg, col_reg}<16'b0001000000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000000000110) && ({row_reg, col_reg}<16'b0001000000001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000000001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001000000001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000000001010) && ({row_reg, col_reg}<16'b0001000000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000000001101) && ({row_reg, col_reg}<16'b0001000000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000000010010) && ({row_reg, col_reg}<16'b0001000000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001000000011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000000011010) && ({row_reg, col_reg}<16'b0001000000100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000000100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000000100010) && ({row_reg, col_reg}<16'b0001000000101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001000000101011) && ({row_reg, col_reg}<16'b0001000000101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001000000101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000000101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000000110000) && ({row_reg, col_reg}<16'b0001000000110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001000000110011) && ({row_reg, col_reg}<16'b0001000000110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000000110110) && ({row_reg, col_reg}<16'b0001000001000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001000001000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000001000001) && ({row_reg, col_reg}<16'b0001000001001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000001001010) && ({row_reg, col_reg}<16'b0001000001001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000001001100) && ({row_reg, col_reg}<16'b0001000001010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001000001010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001000001010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000001010110) && ({row_reg, col_reg}<16'b0001000001011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000001011001) && ({row_reg, col_reg}<16'b0001000001011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000001011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000001011110) && ({row_reg, col_reg}<16'b0001000001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001000001100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000001100010) && ({row_reg, col_reg}<16'b0001000001100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000001100100) && ({row_reg, col_reg}<16'b0001000001100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001000001100110) && ({row_reg, col_reg}<16'b0001000001101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001000001101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000001101001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001000001101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000001101011) && ({row_reg, col_reg}<16'b0001000001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000001110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000001110001) && ({row_reg, col_reg}<16'b0001000001111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000001111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000001111010) && ({row_reg, col_reg}<16'b0001000010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000010000001) && ({row_reg, col_reg}<16'b0001000010010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001000010010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000010010100) && ({row_reg, col_reg}<16'b0001000010010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000010010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000010010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000010011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000010011001) && ({row_reg, col_reg}<16'b0001000010011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001000010011101) && ({row_reg, col_reg}<16'b0001000010100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000010100000) && ({row_reg, col_reg}<16'b0001000010100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000010100010) && ({row_reg, col_reg}<16'b0001000010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000010100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001000010100110) && ({row_reg, col_reg}<16'b0001000010101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001000010101001) && ({row_reg, col_reg}<16'b0001000010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000010101101) && ({row_reg, col_reg}<16'b0001000010101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000010101111) && ({row_reg, col_reg}<16'b0001000010110001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001000010110001) && ({row_reg, col_reg}<16'b0001000010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001000010110101) && ({row_reg, col_reg}<16'b0001000010111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001000010111000) && ({row_reg, col_reg}<16'b0001000010111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001000010111011) && ({row_reg, col_reg}<16'b0001000010111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001000010111101) && ({row_reg, col_reg}<16'b0001000011000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000011000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001000011000010) && ({row_reg, col_reg}<16'b0001000011000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000011000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000011000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000011000110) && ({row_reg, col_reg}<16'b0001000011001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001000011001010) && ({row_reg, col_reg}<16'b0001000011001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000011001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000011001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000011001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000011001111)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0001000011010000) && ({row_reg, col_reg}<16'b0001000011010010)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0001000011010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001000011010011) && ({row_reg, col_reg}<16'b0001000011010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000011010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001000011010111) && ({row_reg, col_reg}<16'b0001000011011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000011011001)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0001000011011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001000011011011) && ({row_reg, col_reg}<16'b0001000011100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001000011100000) && ({row_reg, col_reg}<16'b0001000011100010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001000011100010) && ({row_reg, col_reg}<16'b0001000011101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001000011101000) && ({row_reg, col_reg}<16'b0001000011101011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001000011101011) && ({row_reg, col_reg}<16'b0001000011101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000011101110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001000011101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001000011110000) && ({row_reg, col_reg}<16'b0001000011110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000011110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000011110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000011110100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001000011110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001000011110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000011110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001000011111000) && ({row_reg, col_reg}<16'b0001000011111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000011111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001000011111100) && ({row_reg, col_reg}<16'b0001000011111110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001000011111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0001000011111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001000100000000) && ({row_reg, col_reg}<16'b0001000100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000100000110) && ({row_reg, col_reg}<16'b0001000100001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000100001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000100001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000100001111) && ({row_reg, col_reg}<16'b0001000100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000100010010) && ({row_reg, col_reg}<16'b0001000100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001000100011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000100011010) && ({row_reg, col_reg}<16'b0001000100100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000100100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000100100010) && ({row_reg, col_reg}<16'b0001000100101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001000100101011) && ({row_reg, col_reg}<16'b0001000100101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000100101101) && ({row_reg, col_reg}<16'b0001000100101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000100101111) && ({row_reg, col_reg}<16'b0001000100110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000100110001) && ({row_reg, col_reg}<16'b0001000100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001000100110011) && ({row_reg, col_reg}<16'b0001000100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000100110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000100110110) && ({row_reg, col_reg}<16'b0001000101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001000101000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000101000001) && ({row_reg, col_reg}<16'b0001000101001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000101001010) && ({row_reg, col_reg}<16'b0001000101001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000101001100) && ({row_reg, col_reg}<16'b0001000101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001000101010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000101010100) && ({row_reg, col_reg}<16'b0001000101010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000101010110) && ({row_reg, col_reg}<16'b0001000101011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000101011001) && ({row_reg, col_reg}<16'b0001000101011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000101011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000101011110) && ({row_reg, col_reg}<16'b0001000101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001000101100001) && ({row_reg, col_reg}<16'b0001000101100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000101100100) && ({row_reg, col_reg}<16'b0001000101101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001000101101000) && ({row_reg, col_reg}<16'b0001000101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001000101101010) && ({row_reg, col_reg}<16'b0001000101101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000101101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000101101101) && ({row_reg, col_reg}<16'b0001000101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000101101111) && ({row_reg, col_reg}<16'b0001000101110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001000101110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000101110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000101110011) && ({row_reg, col_reg}<16'b0001000101110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000101110111) && ({row_reg, col_reg}<16'b0001000101111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000101111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000101111010) && ({row_reg, col_reg}<16'b0001000101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000101111111) && ({row_reg, col_reg}<16'b0001000110000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000110000001) && ({row_reg, col_reg}<16'b0001000110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001000110010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000110010101) && ({row_reg, col_reg}<16'b0001000110011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000110011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001000110011001) && ({row_reg, col_reg}<16'b0001000110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001000110011101) && ({row_reg, col_reg}<16'b0001000110100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000110100000) && ({row_reg, col_reg}<16'b0001000110100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001000110100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000110100011) && ({row_reg, col_reg}<16'b0001000110100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000110100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001000110101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000110101010) && ({row_reg, col_reg}<16'b0001000110101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001000110101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000110101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001000110101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001000110101111) && ({row_reg, col_reg}<16'b0001000110110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001000110110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001000110110010) && ({row_reg, col_reg}<16'b0001000110110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001000110110100) && ({row_reg, col_reg}<16'b0001000110111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000110111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001000110111010) && ({row_reg, col_reg}<16'b0001000110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001000110111110) && ({row_reg, col_reg}<16'b0001000111000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000111000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001000111000010) && ({row_reg, col_reg}<16'b0001000111000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001000111000100) && ({row_reg, col_reg}<16'b0001000111000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001000111000110) && ({row_reg, col_reg}<16'b0001000111001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001000111001001) && ({row_reg, col_reg}<16'b0001000111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001000111001011) && ({row_reg, col_reg}<16'b0001000111001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000111001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000111001110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0001000111001111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001000111010000)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0001000111010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001000111010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001000111010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001000111010100) && ({row_reg, col_reg}<16'b0001000111011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001000111011001) && ({row_reg, col_reg}<16'b0001000111011011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001000111011011) && ({row_reg, col_reg}<16'b0001000111011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000111011111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001000111100000) && ({row_reg, col_reg}<16'b0001000111100010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001000111100010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001000111100011) && ({row_reg, col_reg}<16'b0001000111100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000111100110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001000111100111) && ({row_reg, col_reg}<16'b0001000111101010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001000111101010) && ({row_reg, col_reg}<16'b0001000111101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000111101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000111110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001000111110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000111110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000111110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001000111110100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001000111110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001000111110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001000111110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001000111111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001000111111001) && ({row_reg, col_reg}<16'b0001000111111011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001000111111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001000111111100) && ({row_reg, col_reg}<16'b0001000111111110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001000111111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0001000111111111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001001000000000) && ({row_reg, col_reg}<16'b0001001000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001000000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001001000000111) && ({row_reg, col_reg}<16'b0001001000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001001000001001) && ({row_reg, col_reg}<16'b0001001000001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001000001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001000001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001001000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001000010000) && ({row_reg, col_reg}<16'b0001001000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001000010010) && ({row_reg, col_reg}<16'b0001001000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001001000011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001000011010) && ({row_reg, col_reg}<16'b0001001000100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001000100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001000100010) && ({row_reg, col_reg}<16'b0001001000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001001000101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001000101011) && ({row_reg, col_reg}<16'b0001001000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001000110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001001000110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001001000110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001000110011) && ({row_reg, col_reg}<16'b0001001000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001000110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001000110110) && ({row_reg, col_reg}<16'b0001001000111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001001000111100) && ({row_reg, col_reg}<16'b0001001000111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001000111110) && ({row_reg, col_reg}<16'b0001001001000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001001001000001) && ({row_reg, col_reg}<16'b0001001001001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001001001010) && ({row_reg, col_reg}<16'b0001001001001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001001001100) && ({row_reg, col_reg}<16'b0001001001010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001001001010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001001010100) && ({row_reg, col_reg}<16'b0001001001010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001001010111) && ({row_reg, col_reg}<16'b0001001001011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001001011001) && ({row_reg, col_reg}<16'b0001001001011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001001011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001001011110) && ({row_reg, col_reg}<16'b0001001001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001001001100001) && ({row_reg, col_reg}<16'b0001001001100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001001100011) && ({row_reg, col_reg}<16'b0001001001100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001001100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001001100110) && ({row_reg, col_reg}<16'b0001001001101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001001101101) && ({row_reg, col_reg}<16'b0001001001110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001001110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001001110011) && ({row_reg, col_reg}<16'b0001001001111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001001111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001001111010) && ({row_reg, col_reg}<16'b0001001010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001010000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001001010000001) && ({row_reg, col_reg}<16'b0001001010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001001010010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001010010101) && ({row_reg, col_reg}<16'b0001001010011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001010011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001010011010) && ({row_reg, col_reg}<16'b0001001010011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001001010011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001010011101) && ({row_reg, col_reg}<16'b0001001010100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001010100000) && ({row_reg, col_reg}<16'b0001001010100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001001010100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001010100011) && ({row_reg, col_reg}<16'b0001001010100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001001010100101) && ({row_reg, col_reg}<16'b0001001010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001001010101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001010101011) && ({row_reg, col_reg}<16'b0001001010101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001010101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001010101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001001010101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001001010110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001010110001) && ({row_reg, col_reg}<16'b0001001010110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001001010110100) && ({row_reg, col_reg}<16'b0001001010110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001010110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001001010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001010111001) && ({row_reg, col_reg}<16'b0001001010111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001010111011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0001001010111100) && ({row_reg, col_reg}<16'b0001001010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001010111110) && ({row_reg, col_reg}<16'b0001001011000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001011000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001011000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001011000100) && ({row_reg, col_reg}<16'b0001001011000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001011000111) && ({row_reg, col_reg}<16'b0001001011001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001011001001) && ({row_reg, col_reg}<16'b0001001011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001011001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001001011001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001011001101) && ({row_reg, col_reg}<16'b0001001011001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001011001111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001001011010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001011010001)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}==16'b0001001011010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001001011010011) && ({row_reg, col_reg}<16'b0001001011010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001011010101) && ({row_reg, col_reg}<16'b0001001011010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001011010111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001001011011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001011011001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0001001011011010) && ({row_reg, col_reg}<16'b0001001011011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001001011011100) && ({row_reg, col_reg}<16'b0001001011011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001001011011110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001001011011111) && ({row_reg, col_reg}<16'b0001001011100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001001011100100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001001011100101) && ({row_reg, col_reg}<16'b0001001011101000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001001011101000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0001001011101001) && ({row_reg, col_reg}<16'b0001001011101011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001001011101011) && ({row_reg, col_reg}<16'b0001001011101101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0001001011101101) && ({row_reg, col_reg}<16'b0001001011101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001001011101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001001011110000) && ({row_reg, col_reg}<16'b0001001011110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001011110011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001001011110100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001001011110101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001001011110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001011110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001011111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001011111001) && ({row_reg, col_reg}<16'b0001001011111011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001001011111011)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0001001011111100) && ({row_reg, col_reg}<16'b0001001011111110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001001011111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0001001011111111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001001100000000) && ({row_reg, col_reg}<16'b0001001100000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001100000111) && ({row_reg, col_reg}<16'b0001001100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001100001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001100001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001100001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001001100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001100001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001001100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001100010000) && ({row_reg, col_reg}<16'b0001001100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001100010010) && ({row_reg, col_reg}<16'b0001001100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001001100011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001100011010) && ({row_reg, col_reg}<16'b0001001100100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001100100001) && ({row_reg, col_reg}<16'b0001001100100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001100100011) && ({row_reg, col_reg}<16'b0001001100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001001100101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001100101011) && ({row_reg, col_reg}<16'b0001001100110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001100110001) && ({row_reg, col_reg}<16'b0001001100110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001001100110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001100110100) && ({row_reg, col_reg}<16'b0001001100110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001100110110) && ({row_reg, col_reg}<16'b0001001100111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001001100111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001100111001) && ({row_reg, col_reg}<16'b0001001100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001001100111100) && ({row_reg, col_reg}<16'b0001001100111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001100111110) && ({row_reg, col_reg}<16'b0001001101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001001101000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001101000001) && ({row_reg, col_reg}<16'b0001001101001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001101001010) && ({row_reg, col_reg}<16'b0001001101001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001101001100) && ({row_reg, col_reg}<16'b0001001101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001001101010001) && ({row_reg, col_reg}<16'b0001001101010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001101010100) && ({row_reg, col_reg}<16'b0001001101011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001101011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001101011110) && ({row_reg, col_reg}<16'b0001001101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001001101100001) && ({row_reg, col_reg}<16'b0001001101100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001101100100) && ({row_reg, col_reg}<16'b0001001101101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001101101001) && ({row_reg, col_reg}<16'b0001001101101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001101101011) && ({row_reg, col_reg}<16'b0001001101101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001101101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001101110000) && ({row_reg, col_reg}<16'b0001001101110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001101110010) && ({row_reg, col_reg}<16'b0001001101110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001101110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001101110101) && ({row_reg, col_reg}<16'b0001001101110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001101110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001001101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001101111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001001101111010) && ({row_reg, col_reg}<16'b0001001101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001001110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001110000001) && ({row_reg, col_reg}<16'b0001001110010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001001110010101) && ({row_reg, col_reg}<16'b0001001110011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001001110011000) && ({row_reg, col_reg}<16'b0001001110100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001110100000) && ({row_reg, col_reg}<16'b0001001110100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001001110100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001110100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001110100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001001110100110) && ({row_reg, col_reg}<16'b0001001110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001001110101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001001110101011) && ({row_reg, col_reg}<16'b0001001110101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001110101101) && ({row_reg, col_reg}<16'b0001001110101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001110101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001110110000) && ({row_reg, col_reg}<16'b0001001110110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001001110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001110110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001110110101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0001001110110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001110110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001001110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001110111001) && ({row_reg, col_reg}<16'b0001001110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001001110111011) && ({row_reg, col_reg}<16'b0001001110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001110111110) && ({row_reg, col_reg}<16'b0001001111000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001111000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001111000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001001111000100) && ({row_reg, col_reg}<16'b0001001111000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001001111000110) && ({row_reg, col_reg}<16'b0001001111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001001111001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001111001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001111001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001001111001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001001111001101) && ({row_reg, col_reg}<16'b0001001111010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001111010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001111010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001001111010010)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==16'b0001001111010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001001111010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001001111010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001111010110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0001001111010111) && ({row_reg, col_reg}<16'b0001001111011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001001111011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001001111011010) && ({row_reg, col_reg}<16'b0001001111011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001001111011100) && ({row_reg, col_reg}<16'b0001001111011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001001111011111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001001111100000) && ({row_reg, col_reg}<16'b0001001111100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001001111100111) && ({row_reg, col_reg}<16'b0001001111101010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001001111101010)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0001001111101011) && ({row_reg, col_reg}<16'b0001001111101101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0001001111101101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0001001111101110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001001111101111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001001111110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001001111110001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001001111110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001001111110011) && ({row_reg, col_reg}<16'b0001001111110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001001111110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001001111110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001111110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001001111111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001001111111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001001111111010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0001001111111011)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0001001111111100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001001111111101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001001111111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0001001111111111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0001010000000000) && ({row_reg, col_reg}<16'b0001010000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010000000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001010000000111) && ({row_reg, col_reg}<16'b0001010000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001010000001001) && ({row_reg, col_reg}<16'b0001010000001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010000001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001010000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010000001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001010000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010000010000) && ({row_reg, col_reg}<16'b0001010000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010000010010) && ({row_reg, col_reg}<16'b0001010000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001010000011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010000011010) && ({row_reg, col_reg}<16'b0001010000100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010000100001) && ({row_reg, col_reg}<16'b0001010000100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010000100011) && ({row_reg, col_reg}<16'b0001010000101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001010000101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010000101100) && ({row_reg, col_reg}<16'b0001010000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010000110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010000110010) && ({row_reg, col_reg}<16'b0001010000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010000110100) && ({row_reg, col_reg}<16'b0001010000110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010000110110) && ({row_reg, col_reg}<16'b0001010001000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001010001000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010001000001) && ({row_reg, col_reg}<16'b0001010001001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010001001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010001001011) && ({row_reg, col_reg}<16'b0001010001010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001010001010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010001010100) && ({row_reg, col_reg}<16'b0001010001011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010001011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010001011110) && ({row_reg, col_reg}<16'b0001010001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001010001100001) && ({row_reg, col_reg}<16'b0001010001100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010001100100) && ({row_reg, col_reg}<16'b0001010001101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010001101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001010001101001) && ({row_reg, col_reg}<16'b0001010001101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010001101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010001101100) && ({row_reg, col_reg}<16'b0001010001110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010001110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001010001110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010001110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010001110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010001110110) && ({row_reg, col_reg}<16'b0001010001111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001010001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010001111001) && ({row_reg, col_reg}<16'b0001010001111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010001111011) && ({row_reg, col_reg}<16'b0001010010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010010000001) && ({row_reg, col_reg}<16'b0001010010010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001010010010101) && ({row_reg, col_reg}<16'b0001010010011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001010010011000) && ({row_reg, col_reg}<16'b0001010010011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010010011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001010010011011) && ({row_reg, col_reg}<16'b0001010010100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010010100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001010010100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001010010100010) && ({row_reg, col_reg}<16'b0001010010100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010010100110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001010010100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001010010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001010010101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001010010101010) && ({row_reg, col_reg}<16'b0001010010101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010010101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010010101110) && ({row_reg, col_reg}<16'b0001010010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010010110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001010010110001) && ({row_reg, col_reg}<16'b0001010010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010010110011) && ({row_reg, col_reg}<16'b0001010010110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010010110110) && ({row_reg, col_reg}<16'b0001010010111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001010010111000) && ({row_reg, col_reg}<16'b0001010010111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001010010111011) && ({row_reg, col_reg}<16'b0001010010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010010111110) && ({row_reg, col_reg}<16'b0001010011000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010011000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010011000100) && ({row_reg, col_reg}<16'b0001010011000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001010011000110) && ({row_reg, col_reg}<16'b0001010011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010011001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010011001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001010011001011) && ({row_reg, col_reg}<16'b0001010011001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010011001101) && ({row_reg, col_reg}<16'b0001010011010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010011010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010011010001) && ({row_reg, col_reg}<16'b0001010011010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001010011010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010011010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001010011010101) && ({row_reg, col_reg}<16'b0001010011010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010011010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001010011011000) && ({row_reg, col_reg}<16'b0001010011011010)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0001010011011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001010011011011) && ({row_reg, col_reg}<16'b0001010011011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010011011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001010011011111) && ({row_reg, col_reg}<16'b0001010011100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001010011100001) && ({row_reg, col_reg}<16'b0001010011100011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001010011100011) && ({row_reg, col_reg}<16'b0001010011100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010011100101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001010011100110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001010011100111) && ({row_reg, col_reg}<16'b0001010011101001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001010011101001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0001010011101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001010011101011) && ({row_reg, col_reg}<16'b0001010011101101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0001010011101101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0001010011101110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001010011101111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001010011110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001010011110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010011110010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001010011110011) && ({row_reg, col_reg}<16'b0001010011110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010011110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010011110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010011110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010011111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010011111001) && ({row_reg, col_reg}<16'b0001010011111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010011111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001010011111100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010011111101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001010011111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0001010011111111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0001010100000000) && ({row_reg, col_reg}<16'b0001010100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010100000110) && ({row_reg, col_reg}<16'b0001010100001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001010100001011) && ({row_reg, col_reg}<16'b0001010100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010100001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001010100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010100010000) && ({row_reg, col_reg}<16'b0001010100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010100010010) && ({row_reg, col_reg}<16'b0001010100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001010100011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010100011010) && ({row_reg, col_reg}<16'b0001010100100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010100100001) && ({row_reg, col_reg}<16'b0001010100100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010100100011) && ({row_reg, col_reg}<16'b0001010100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001010100101010) && ({row_reg, col_reg}<16'b0001010100101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010100101100) && ({row_reg, col_reg}<16'b0001010100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010100110100) && ({row_reg, col_reg}<16'b0001010100110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010100110110) && ({row_reg, col_reg}<16'b0001010101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001010101000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010101000001) && ({row_reg, col_reg}<16'b0001010101001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010101001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010101001011) && ({row_reg, col_reg}<16'b0001010101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001010101010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010101010100) && ({row_reg, col_reg}<16'b0001010101011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010101011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010101011110) && ({row_reg, col_reg}<16'b0001010101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001010101100001) && ({row_reg, col_reg}<16'b0001010101100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010101100011) && ({row_reg, col_reg}<16'b0001010101100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010101100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010101100110) && ({row_reg, col_reg}<16'b0001010101101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010101101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010101101001) && ({row_reg, col_reg}<16'b0001010101101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001010101101011) && ({row_reg, col_reg}<16'b0001010101101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010101101101) && ({row_reg, col_reg}<16'b0001010101101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010101101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001010101110000) && ({row_reg, col_reg}<16'b0001010101110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010101110010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0001010101110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010101110100) && ({row_reg, col_reg}<16'b0001010101110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001010101110110) && ({row_reg, col_reg}<16'b0001010101111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010101111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001010101111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001010101111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001010101111100) && ({row_reg, col_reg}<16'b0001010110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010110000001) && ({row_reg, col_reg}<16'b0001010110010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001010110010101) && ({row_reg, col_reg}<16'b0001010110011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001010110011011) && ({row_reg, col_reg}<16'b0001010110100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010110100000) && ({row_reg, col_reg}<16'b0001010110100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001010110100011) && ({row_reg, col_reg}<16'b0001010110100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001010110100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001010110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001010110101001) && ({row_reg, col_reg}<16'b0001010110101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001010110101110) && ({row_reg, col_reg}<16'b0001010110110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001010110110001) && ({row_reg, col_reg}<16'b0001010110110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001010110110011) && ({row_reg, col_reg}<16'b0001010110110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010110110110) && ({row_reg, col_reg}<16'b0001010110111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001010110111000) && ({row_reg, col_reg}<16'b0001010110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010110111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010110111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010110111101) && ({row_reg, col_reg}<16'b0001010111000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010111000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010111000011) && ({row_reg, col_reg}<16'b0001010111000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010111000101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001010111000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010111001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001010111001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001010111001010) && ({row_reg, col_reg}<16'b0001010111001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001010111001101) && ({row_reg, col_reg}<16'b0001010111001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010111001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010111010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010111010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001010111010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001010111010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001010111010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010111010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010111010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001010111010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010111011000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001010111011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001010111011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001010111011011) && ({row_reg, col_reg}<16'b0001010111011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010111011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001010111011111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001010111100000) && ({row_reg, col_reg}<16'b0001010111100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010111100010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001010111100011) && ({row_reg, col_reg}<16'b0001010111100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010111100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001010111100110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010111100111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0001010111101000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0001010111101001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010111101010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001010111101011) && ({row_reg, col_reg}<16'b0001010111101101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0001010111101101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0001010111101110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001010111101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010111110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010111110001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001010111110010) && ({row_reg, col_reg}<16'b0001010111110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010111110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010111110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010111110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001010111111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001010111111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001010111111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001010111111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001010111111100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001010111111101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001010111111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0001010111111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011000000000) && ({row_reg, col_reg}<16'b0001011000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011000000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011000000110) && ({row_reg, col_reg}<16'b0001011000001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001011000001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001011000001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011000001100) && ({row_reg, col_reg}<16'b0001011000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011000010000) && ({row_reg, col_reg}<16'b0001011000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011000010010) && ({row_reg, col_reg}<16'b0001011000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001011000011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011000011010) && ({row_reg, col_reg}<16'b0001011000100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011000100001) && ({row_reg, col_reg}<16'b0001011000100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011000100011) && ({row_reg, col_reg}<16'b0001011000101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001011000101001) && ({row_reg, col_reg}<16'b0001011000101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011000101011) && ({row_reg, col_reg}<16'b0001011000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011000110100) && ({row_reg, col_reg}<16'b0001011000110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011000110110) && ({row_reg, col_reg}<16'b0001011001000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001011001000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011001000001) && ({row_reg, col_reg}<16'b0001011001001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011001001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011001001010) && ({row_reg, col_reg}<16'b0001011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001011001010001) && ({row_reg, col_reg}<16'b0001011001010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011001010100) && ({row_reg, col_reg}<16'b0001011001011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011001011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011001011110) && ({row_reg, col_reg}<16'b0001011001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001011001100001) && ({row_reg, col_reg}<16'b0001011001100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011001100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001011001100100) && ({row_reg, col_reg}<16'b0001011001100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011001100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001011001101000) && ({row_reg, col_reg}<16'b0001011001101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011001101010) && ({row_reg, col_reg}<16'b0001011001101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001011001101111) && ({row_reg, col_reg}<16'b0001011001110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011001110001) && ({row_reg, col_reg}<16'b0001011001110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001011001110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011001110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001011001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011001111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011001111010) && ({row_reg, col_reg}<16'b0001011001111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001011001111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011001111101) && ({row_reg, col_reg}<16'b0001011010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011010000010) && ({row_reg, col_reg}<16'b0001011010010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001011010010101) && ({row_reg, col_reg}<16'b0001011010011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001011010011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011010011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011010011101) && ({row_reg, col_reg}<16'b0001011010100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011010100000) && ({row_reg, col_reg}<16'b0001011010100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001011010100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001011010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001011010100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011010101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001011010101001) && ({row_reg, col_reg}<16'b0001011010101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011010101110) && ({row_reg, col_reg}<16'b0001011010110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001011010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011010110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011010110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001011010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011010110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001011010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011010111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011010111011) && ({row_reg, col_reg}<16'b0001011010111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001011010111101) && ({row_reg, col_reg}<16'b0001011010111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011010111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001011011000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011011000001) && ({row_reg, col_reg}<16'b0001011011000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011011000011) && ({row_reg, col_reg}<16'b0001011011000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011011000101) && ({row_reg, col_reg}<16'b0001011011000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011011000111) && ({row_reg, col_reg}<16'b0001011011001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001011011001001) && ({row_reg, col_reg}<16'b0001011011001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011011001110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0001011011001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001011011010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011011010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011011010010) && ({row_reg, col_reg}<16'b0001011011010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001011011010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011011010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011011010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011011010111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001011011011000) && ({row_reg, col_reg}<16'b0001011011011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011011011010) && ({row_reg, col_reg}<16'b0001011011011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001011011011100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0001011011011101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001011011011110) && ({row_reg, col_reg}<16'b0001011011100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011011100010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001011011100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001011011100100) && ({row_reg, col_reg}<16'b0001011011100111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001011011100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001011011101000) && ({row_reg, col_reg}<16'b0001011011101010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001011011101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001011011101011)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0001011011101100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0001011011101101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0001011011101110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0001011011101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0001011011110000) && ({row_reg, col_reg}<16'b0001011011110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001011011110010) && ({row_reg, col_reg}<16'b0001011011110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001011011110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011011110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011011110111) && ({row_reg, col_reg}<16'b0001011011111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011011111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001011011111010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0001011011111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001011011111100) && ({row_reg, col_reg}<16'b0001011011111110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001011011111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0001011011111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011100000000) && ({row_reg, col_reg}<16'b0001011100000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011100000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001011100000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011100000101) && ({row_reg, col_reg}<16'b0001011100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011100000111) && ({row_reg, col_reg}<16'b0001011100001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011100001001) && ({row_reg, col_reg}<16'b0001011100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011100001100) && ({row_reg, col_reg}<16'b0001011100001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011100001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011100001111) && ({row_reg, col_reg}<16'b0001011100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011100010010) && ({row_reg, col_reg}<16'b0001011100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001011100011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011100011010) && ({row_reg, col_reg}<16'b0001011100100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011100100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011100100011) && ({row_reg, col_reg}<16'b0001011100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001011100101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011100101011) && ({row_reg, col_reg}<16'b0001011100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011100110100) && ({row_reg, col_reg}<16'b0001011100110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011100110110) && ({row_reg, col_reg}<16'b0001011101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001011101000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011101000001) && ({row_reg, col_reg}<16'b0001011101001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011101001001) && ({row_reg, col_reg}<16'b0001011101001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011101001011) && ({row_reg, col_reg}<16'b0001011101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001011101010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011101010100) && ({row_reg, col_reg}<16'b0001011101011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011101011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011101011110) && ({row_reg, col_reg}<16'b0001011101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001011101100001) && ({row_reg, col_reg}<16'b0001011101100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011101100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001011101100100) && ({row_reg, col_reg}<16'b0001011101100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011101100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001011101101000) && ({row_reg, col_reg}<16'b0001011101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011101101010) && ({row_reg, col_reg}<16'b0001011101101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001011101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011101110000) && ({row_reg, col_reg}<16'b0001011101110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011101110010) && ({row_reg, col_reg}<16'b0001011101110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001011101110110) && ({row_reg, col_reg}<16'b0001011101111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011101111000) && ({row_reg, col_reg}<16'b0001011101111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011101111100) && ({row_reg, col_reg}<16'b0001011101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011101111110) && ({row_reg, col_reg}<16'b0001011110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011110000001) && ({row_reg, col_reg}<16'b0001011110010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001011110010101) && ({row_reg, col_reg}<16'b0001011110011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011110011011) && ({row_reg, col_reg}<16'b0001011110011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001011110011101) && ({row_reg, col_reg}<16'b0001011110100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011110100000) && ({row_reg, col_reg}<16'b0001011110100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001011110100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001011110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011110100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001011110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001011110101001) && ({row_reg, col_reg}<16'b0001011110101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001011110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011110101110) && ({row_reg, col_reg}<16'b0001011110110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001011110110011) && ({row_reg, col_reg}<16'b0001011110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011110110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001011110110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011110110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001011110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001011110111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011110111011) && ({row_reg, col_reg}<16'b0001011110111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001011110111101) && ({row_reg, col_reg}<16'b0001011110111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011110111111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001011111000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011111000001) && ({row_reg, col_reg}<16'b0001011111000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011111000011) && ({row_reg, col_reg}<16'b0001011111001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001011111001000) && ({row_reg, col_reg}<16'b0001011111001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011111001010) && ({row_reg, col_reg}<16'b0001011111001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011111001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001011111001110) && ({row_reg, col_reg}<16'b0001011111010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001011111010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001011111010001) && ({row_reg, col_reg}<16'b0001011111010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001011111010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011111010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011111010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001011111010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011111011000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0001011111011001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0001011111011010) && ({row_reg, col_reg}<16'b0001011111011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001011111011100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0001011111011101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001011111011110) && ({row_reg, col_reg}<16'b0001011111100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011111100000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001011111100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001011111100010) && ({row_reg, col_reg}<16'b0001011111100100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001011111100100) && ({row_reg, col_reg}<16'b0001011111101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011111101000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001011111101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011111101010)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0001011111101011) && ({row_reg, col_reg}<16'b0001011111101101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0001011111101101) && ({row_reg, col_reg}<16'b0001011111101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001011111101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001011111110000) && ({row_reg, col_reg}<16'b0001011111110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001011111110010) && ({row_reg, col_reg}<16'b0001011111110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001011111110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001011111110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001011111110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011111111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001011111111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001011111111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001011111111011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0001011111111100) && ({row_reg, col_reg}<16'b0001011111111110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001011111111110)) color_data = 12'b010000110001;

		if(({row_reg, col_reg}==16'b0001011111111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100000000000) && ({row_reg, col_reg}<16'b0001100000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100000000101) && ({row_reg, col_reg}<16'b0001100000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001100000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100000001101) && ({row_reg, col_reg}<16'b0001100000001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100000001111) && ({row_reg, col_reg}<16'b0001100000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100000010010) && ({row_reg, col_reg}<16'b0001100000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001100000011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100000011010) && ({row_reg, col_reg}<16'b0001100000100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100000100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100000100100) && ({row_reg, col_reg}<16'b0001100000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001100000101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100000101011) && ({row_reg, col_reg}<16'b0001100000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100000110100) && ({row_reg, col_reg}<16'b0001100000110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100000110110) && ({row_reg, col_reg}<16'b0001100001000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001100001000001) && ({row_reg, col_reg}<16'b0001100001001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100001001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100001001100) && ({row_reg, col_reg}<16'b0001100001010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001100001010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100001010100) && ({row_reg, col_reg}<16'b0001100001011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100001011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100001011110) && ({row_reg, col_reg}<16'b0001100001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001100001100001) && ({row_reg, col_reg}<16'b0001100001100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100001100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001100001100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100001100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001100001100110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001100001100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001100001101000) && ({row_reg, col_reg}<16'b0001100001101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100001101010) && ({row_reg, col_reg}<16'b0001100001110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001100001110011) && ({row_reg, col_reg}<16'b0001100001110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100001110101) && ({row_reg, col_reg}<16'b0001100001110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001100001110111) && ({row_reg, col_reg}<16'b0001100001111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001100001111010) && ({row_reg, col_reg}<16'b0001100001111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100001111100) && ({row_reg, col_reg}<16'b0001100010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100010000001) && ({row_reg, col_reg}<16'b0001100010010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001100010010101) && ({row_reg, col_reg}<16'b0001100010011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100010011011) && ({row_reg, col_reg}<16'b0001100010011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001100010011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100010011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001100010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100010100000) && ({row_reg, col_reg}<16'b0001100010100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001100010100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001100010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100010100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001100010100110) && ({row_reg, col_reg}<16'b0001100010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001100010101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100010101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001100010101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100010101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001100010101101) && ({row_reg, col_reg}<16'b0001100010101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100010101111) && ({row_reg, col_reg}<16'b0001100010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001100010110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001100010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100010110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001100010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001100010110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001100010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100010111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100010111011) && ({row_reg, col_reg}<16'b0001100010111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001100010111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100010111110) && ({row_reg, col_reg}<16'b0001100011000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100011000010) && ({row_reg, col_reg}<16'b0001100011000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100011000100) && ({row_reg, col_reg}<16'b0001100011001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100011001011) && ({row_reg, col_reg}<16'b0001100011001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001100011001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100011001110) && ({row_reg, col_reg}<16'b0001100011010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001100011010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100011010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100011010010) && ({row_reg, col_reg}<16'b0001100011010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001100011010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100011010101) && ({row_reg, col_reg}<16'b0001100011010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100011010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001100011011000) && ({row_reg, col_reg}<16'b0001100011011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001100011011100) && ({row_reg, col_reg}<16'b0001100011011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100011011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001100011011111) && ({row_reg, col_reg}<16'b0001100011100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100011100010) && ({row_reg, col_reg}<16'b0001100011100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001100011100101) && ({row_reg, col_reg}<16'b0001100011101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100011101001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001100011101010) && ({row_reg, col_reg}<16'b0001100011110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100011110010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001100011110011) && ({row_reg, col_reg}<16'b0001100011110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001100011110101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001100011110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100011110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001100011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001100011111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100011111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001100011111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100011111100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001100011111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100011111110)) color_data = 12'b010000100001;

		if(({row_reg, col_reg}==16'b0001100011111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100100000000) && ({row_reg, col_reg}<16'b0001100100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100100000101) && ({row_reg, col_reg}<16'b0001100100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100100001100) && ({row_reg, col_reg}<16'b0001100100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100100010010) && ({row_reg, col_reg}<16'b0001100100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001100100011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100100011010) && ({row_reg, col_reg}<16'b0001100100100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100100100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100100100100) && ({row_reg, col_reg}<16'b0001100100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001100100101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100100101011) && ({row_reg, col_reg}<16'b0001100100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100100110100) && ({row_reg, col_reg}<16'b0001100100110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100100110110) && ({row_reg, col_reg}<16'b0001100101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001100101000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100101000001) && ({row_reg, col_reg}<16'b0001100101001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100101001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100101001100) && ({row_reg, col_reg}<16'b0001100101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001100101010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100101010100) && ({row_reg, col_reg}<16'b0001100101011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100101011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100101011110) && ({row_reg, col_reg}<16'b0001100101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001100101100001) && ({row_reg, col_reg}<16'b0001100101100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100101100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001100101100101) && ({row_reg, col_reg}<16'b0001100101100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001100101100111) && ({row_reg, col_reg}<16'b0001100101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100101101010) && ({row_reg, col_reg}<16'b0001100101101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001100101101100) && ({row_reg, col_reg}<16'b0001100101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100101110000) && ({row_reg, col_reg}<16'b0001100101110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001100101110010) && ({row_reg, col_reg}<16'b0001100101110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100101110101) && ({row_reg, col_reg}<16'b0001100101111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001100101111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001100101111001) && ({row_reg, col_reg}<16'b0001100101111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001100101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100110000001) && ({row_reg, col_reg}<16'b0001100110010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001100110010101) && ({row_reg, col_reg}<16'b0001100110010111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001100110010111) && ({row_reg, col_reg}<16'b0001100110011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100110011010) && ({row_reg, col_reg}<16'b0001100110011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001100110011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100110011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001100110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001100110100000) && ({row_reg, col_reg}<16'b0001100110100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001100110100011) && ({row_reg, col_reg}<16'b0001100110100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100110100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001100110100110) && ({row_reg, col_reg}<16'b0001100110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100110101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001100110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100110101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001100110101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100110101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100110101101) && ({row_reg, col_reg}<16'b0001100110110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001100110110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001100110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100110110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001100110110110) && ({row_reg, col_reg}<16'b0001100110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001100110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100110111001) && ({row_reg, col_reg}<16'b0001100110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100110111011) && ({row_reg, col_reg}<16'b0001100110111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001100110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001100110111110) && ({row_reg, col_reg}<16'b0001100111000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100111000001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001100111000010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001100111000011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0001100111000100) && ({row_reg, col_reg}<16'b0001100111001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100111001000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001100111001001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001100111001010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100111001011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001100111001100)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0001100111001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100111001110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0001100111001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100111010000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001100111010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001100111010010) && ({row_reg, col_reg}<16'b0001100111010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001100111010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001100111010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100111010110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001100111010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100111011000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0001100111011001) && ({row_reg, col_reg}<16'b0001100111011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001100111011101) && ({row_reg, col_reg}<16'b0001100111011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001100111011111) && ({row_reg, col_reg}<16'b0001100111100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001100111100001) && ({row_reg, col_reg}<16'b0001100111100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001100111100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001100111100100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001100111100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100111100110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001100111100111) && ({row_reg, col_reg}<16'b0001100111101010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100111101010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001100111101011) && ({row_reg, col_reg}<16'b0001100111101101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001100111101101) && ({row_reg, col_reg}<16'b0001100111110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100111110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001100111110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100111110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100111110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001100111110100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0001100111110101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001100111110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001100111110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001100111111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001100111111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001100111111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001100111111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001100111111100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001100111111101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001100111111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0001100111111111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001101000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101000000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001101000000010) && ({row_reg, col_reg}<16'b0001101000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101000000101) && ({row_reg, col_reg}<16'b0001101000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001101000001100) && ({row_reg, col_reg}<16'b0001101000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101000010010) && ({row_reg, col_reg}<16'b0001101000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001101000011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101000011010) && ({row_reg, col_reg}<16'b0001101000100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101000100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101000100100) && ({row_reg, col_reg}<16'b0001101000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001101000101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101000101011) && ({row_reg, col_reg}<16'b0001101000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101000110100) && ({row_reg, col_reg}<16'b0001101000110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101000110110) && ({row_reg, col_reg}<16'b0001101001000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001101001000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101001000001) && ({row_reg, col_reg}<16'b0001101001001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101001001010) && ({row_reg, col_reg}<16'b0001101001001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101001001100) && ({row_reg, col_reg}<16'b0001101001010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001101001010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101001010100) && ({row_reg, col_reg}<16'b0001101001011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101001011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101001011110) && ({row_reg, col_reg}<16'b0001101001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001101001100001) && ({row_reg, col_reg}<16'b0001101001100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101001100100) && ({row_reg, col_reg}<16'b0001101001100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001101001100110) && ({row_reg, col_reg}<16'b0001101001101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101001101001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001101001101010) && ({row_reg, col_reg}<16'b0001101001110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001101001110010) && ({row_reg, col_reg}<16'b0001101001110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101001110101) && ({row_reg, col_reg}<16'b0001101001110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001101001110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101001111000) && ({row_reg, col_reg}<16'b0001101001111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101001111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001101001111101) && ({row_reg, col_reg}<16'b0001101010000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001101010000001) && ({row_reg, col_reg}<16'b0001101010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001101010010100) && ({row_reg, col_reg}<16'b0001101010010111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001101010010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101010011000) && ({row_reg, col_reg}<16'b0001101010011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101010011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101010011011) && ({row_reg, col_reg}<16'b0001101010011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101010011101) && ({row_reg, col_reg}<16'b0001101010100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101010100000) && ({row_reg, col_reg}<16'b0001101010100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001101010100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001101010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101010100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001101010100110) && ({row_reg, col_reg}<16'b0001101010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101010101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101010101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101010101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001101010101011) && ({row_reg, col_reg}<16'b0001101010101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001101010101101) && ({row_reg, col_reg}<16'b0001101010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101010110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001101010110011) && ({row_reg, col_reg}<16'b0001101010110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101010110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001101010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001101010111001) && ({row_reg, col_reg}<16'b0001101010111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001101010111011) && ({row_reg, col_reg}<16'b0001101010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001101010111110) && ({row_reg, col_reg}<16'b0001101011000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101011000001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001101011000010)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0001101011000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001101011000100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0001101011000101) && ({row_reg, col_reg}<16'b0001101011001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101011001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001101011001001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001101011001010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101011001011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001101011001100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001101011001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001101011001110) && ({row_reg, col_reg}<16'b0001101011010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001101011010000) && ({row_reg, col_reg}<16'b0001101011010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101011010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101011010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101011010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001101011010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101011010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101011010111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001101011011000) && ({row_reg, col_reg}<16'b0001101011011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001101011011010) && ({row_reg, col_reg}<16'b0001101011011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001101011011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101011011110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001101011011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101011100000) && ({row_reg, col_reg}<16'b0001101011100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001101011100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101011100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101011100100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001101011100101) && ({row_reg, col_reg}<16'b0001101011101011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101011101011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001101011101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101011101101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001101011101110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001101011101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101011110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0001101011110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101011110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001101011110011) && ({row_reg, col_reg}<16'b0001101011110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001101011110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001101011110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101011110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101011111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001101011111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101011111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001101011111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101011111100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001101011111101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001101011111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0001101011111111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0001101100000000) && ({row_reg, col_reg}<16'b0001101100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101100000101) && ({row_reg, col_reg}<16'b0001101100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001101100001100) && ({row_reg, col_reg}<16'b0001101100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101100010010) && ({row_reg, col_reg}<16'b0001101100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001101100011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101100011010) && ({row_reg, col_reg}<16'b0001101100100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101100100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101100100100) && ({row_reg, col_reg}<16'b0001101100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001101100101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101100101011) && ({row_reg, col_reg}<16'b0001101100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101100110100) && ({row_reg, col_reg}<16'b0001101100110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101100110110) && ({row_reg, col_reg}<16'b0001101101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001101101000001) && ({row_reg, col_reg}<16'b0001101101001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101101001010) && ({row_reg, col_reg}<16'b0001101101001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101101001100) && ({row_reg, col_reg}<16'b0001101101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001101101010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101101010100) && ({row_reg, col_reg}<16'b0001101101011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101101011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101101011110) && ({row_reg, col_reg}<16'b0001101101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001101101100001) && ({row_reg, col_reg}<16'b0001101101100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101101100100) && ({row_reg, col_reg}<16'b0001101101100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001101101100110) && ({row_reg, col_reg}<16'b0001101101101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101101101001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001101101101010) && ({row_reg, col_reg}<16'b0001101101110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001101101110001) && ({row_reg, col_reg}<16'b0001101101110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101101110101) && ({row_reg, col_reg}<16'b0001101101110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001101101110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001101101111000) && ({row_reg, col_reg}<16'b0001101101111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001101101111010) && ({row_reg, col_reg}<16'b0001101101111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101101111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001101101111110) && ({row_reg, col_reg}<16'b0001101110000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101110000010) && ({row_reg, col_reg}<16'b0001101110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001101110010100) && ({row_reg, col_reg}<16'b0001101110010110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101110010110) && ({row_reg, col_reg}<16'b0001101110011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101110011000) && ({row_reg, col_reg}<16'b0001101110011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101110011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101110011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101110011100) && ({row_reg, col_reg}<16'b0001101110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101110011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101110100000) && ({row_reg, col_reg}<16'b0001101110100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001101110100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001101110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101110100101) && ({row_reg, col_reg}<16'b0001101110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101110101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001101110101010) && ({row_reg, col_reg}<16'b0001101110101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001101110101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001101110101101) && ({row_reg, col_reg}<16'b0001101110110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101110110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001101110110011) && ({row_reg, col_reg}<16'b0001101110110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101110110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101110110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001101110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001101110111001) && ({row_reg, col_reg}<16'b0001101110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001101110111011) && ({row_reg, col_reg}<16'b0001101110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001101110111101) && ({row_reg, col_reg}<16'b0001101111000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101111000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101111000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001101111000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001101111000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001101111000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101111000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001101111000111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001101111001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001101111001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001101111001010) && ({row_reg, col_reg}<16'b0001101111001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101111001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001101111001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101111010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101111010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001101111010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001101111010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101111010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101111010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101111010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101111010111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001101111011000) && ({row_reg, col_reg}<16'b0001101111011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001101111011010) && ({row_reg, col_reg}<16'b0001101111011110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001101111011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001101111011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001101111100000) && ({row_reg, col_reg}<16'b0001101111100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001101111100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101111100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101111100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001101111100101) && ({row_reg, col_reg}<16'b0001101111100111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001101111100111) && ({row_reg, col_reg}<16'b0001101111101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101111101100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001101111101101) && ({row_reg, col_reg}<16'b0001101111101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001101111101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001101111110000) && ({row_reg, col_reg}<16'b0001101111110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101111110011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001101111110100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001101111110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101111110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001101111110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101111111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001101111111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001101111111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001101111111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001101111111100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001101111111101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001101111111110)) color_data = 12'b010000110001;

		if(({row_reg, col_reg}==16'b0001101111111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001110000000000) && ({row_reg, col_reg}<16'b0001110000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110000000110) && ({row_reg, col_reg}<16'b0001110000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001110000001100) && ({row_reg, col_reg}<16'b0001110000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110000010010) && ({row_reg, col_reg}<16'b0001110000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001110000011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110000011010) && ({row_reg, col_reg}<16'b0001110000100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110000100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110000100100) && ({row_reg, col_reg}<16'b0001110000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001110000101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110000101011) && ({row_reg, col_reg}<16'b0001110000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110000110100) && ({row_reg, col_reg}<16'b0001110000110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110000110110) && ({row_reg, col_reg}<16'b0001110001000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001110001000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110001000001) && ({row_reg, col_reg}<16'b0001110001001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110001001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110001001100) && ({row_reg, col_reg}<16'b0001110001010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001110001010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110001010100) && ({row_reg, col_reg}<16'b0001110001011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110001011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110001011110) && ({row_reg, col_reg}<16'b0001110001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001110001100001) && ({row_reg, col_reg}<16'b0001110001100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110001100100) && ({row_reg, col_reg}<16'b0001110001100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001110001100111) && ({row_reg, col_reg}<16'b0001110001101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110001101001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110001101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001110001101011) && ({row_reg, col_reg}<16'b0001110001101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110001101101) && ({row_reg, col_reg}<16'b0001110001110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001110001110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110001111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001110001111001) && ({row_reg, col_reg}<16'b0001110001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110001111101) && ({row_reg, col_reg}<16'b0001110001111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001110001111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001110010000000) && ({row_reg, col_reg}<16'b0001110010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110010000010) && ({row_reg, col_reg}<16'b0001110010010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001110010010011) && ({row_reg, col_reg}<16'b0001110010010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110010010101) && ({row_reg, col_reg}<16'b0001110010011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110010011000) && ({row_reg, col_reg}<16'b0001110010011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001110010011010) && ({row_reg, col_reg}<16'b0001110010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110010011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110010100000) && ({row_reg, col_reg}<16'b0001110010100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001110010100011) && ({row_reg, col_reg}<16'b0001110010100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110010100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001110010100110) && ({row_reg, col_reg}<16'b0001110010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110010101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001110010101001) && ({row_reg, col_reg}<16'b0001110010101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110010101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001110010101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001110010101101) && ({row_reg, col_reg}<16'b0001110010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110010110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001110010110011) && ({row_reg, col_reg}<16'b0001110010110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110010110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110010111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110010111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110010111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110010111101) && ({row_reg, col_reg}<16'b0001110011000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001110011000001) && ({row_reg, col_reg}<16'b0001110011000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110011000011) && ({row_reg, col_reg}<16'b0001110011000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001110011000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110011000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001110011000111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0001110011001000) && ({row_reg, col_reg}<16'b0001110011001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110011001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001110011001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110011010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110011010001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110011010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110011010011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110011010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110011010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001110011010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110011010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001110011011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110011011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110011011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001110011011011) && ({row_reg, col_reg}<16'b0001110011011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110011011101)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0001110011011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110011011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001110011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001110011100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0001110011100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001110011100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001110011100100) && ({row_reg, col_reg}<16'b0001110011100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110011100110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001110011100111) && ({row_reg, col_reg}<16'b0001110011101011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110011101011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001110011101100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001110011101101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0001110011101110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001110011101111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001110011110000) && ({row_reg, col_reg}<16'b0001110011110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001110011110011) && ({row_reg, col_reg}<16'b0001110011110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001110011110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110011110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001110011110111) && ({row_reg, col_reg}<16'b0001110011111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110011111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110011111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110011111100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001110011111101)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}>=16'b0001110011111110) && ({row_reg, col_reg}<16'b0001110100000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001110100000000) && ({row_reg, col_reg}<16'b0001110100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001110100000010) && ({row_reg, col_reg}<16'b0001110100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110100000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001110100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110100000111) && ({row_reg, col_reg}<16'b0001110100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001110100001100) && ({row_reg, col_reg}<16'b0001110100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110100010010) && ({row_reg, col_reg}<16'b0001110100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001110100011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110100011010) && ({row_reg, col_reg}<16'b0001110100100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110100100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110100100100) && ({row_reg, col_reg}<16'b0001110100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001110100101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110100101011) && ({row_reg, col_reg}<16'b0001110100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110100110100) && ({row_reg, col_reg}<16'b0001110100110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110100110110) && ({row_reg, col_reg}<16'b0001110101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001110101000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110101000001) && ({row_reg, col_reg}<16'b0001110101001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110101001100) && ({row_reg, col_reg}<16'b0001110101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001110101010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110101010100) && ({row_reg, col_reg}<16'b0001110101011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110101011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110101011110) && ({row_reg, col_reg}<16'b0001110101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001110101100001) && ({row_reg, col_reg}<16'b0001110101100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110101100100) && ({row_reg, col_reg}<16'b0001110101101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001110101101000) && ({row_reg, col_reg}<16'b0001110101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110101101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001110101101011) && ({row_reg, col_reg}<16'b0001110101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110101101110) && ({row_reg, col_reg}<16'b0001110101110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001110101110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110101110100) && ({row_reg, col_reg}<16'b0001110101110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001110101110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110101111000) && ({row_reg, col_reg}<16'b0001110101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001110101111011) && ({row_reg, col_reg}<16'b0001110101111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110101111101) && ({row_reg, col_reg}<16'b0001110101111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001110101111111) && ({row_reg, col_reg}<16'b0001110110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110110000010) && ({row_reg, col_reg}<16'b0001110110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001110110010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110110010101) && ({row_reg, col_reg}<16'b0001110110011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110110011000) && ({row_reg, col_reg}<16'b0001110110011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001110110011010) && ({row_reg, col_reg}<16'b0001110110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110110011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110110100000) && ({row_reg, col_reg}<16'b0001110110100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001110110100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001110110100011) && ({row_reg, col_reg}<16'b0001110110100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110110100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001110110100110) && ({row_reg, col_reg}<16'b0001110110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110110101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001110110101010) && ({row_reg, col_reg}<16'b0001110110110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110110110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110110110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110110110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110110110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110110111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110110111010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0001110110111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001110110111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110110111110) && ({row_reg, col_reg}<16'b0001110111000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001110111000010) && ({row_reg, col_reg}<16'b0001110111001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110111001010) && ({row_reg, col_reg}<16'b0001110111001100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110111001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001110111001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110111001110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110111001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110111010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001110111010001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110111010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001110111010011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001110111010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110111010101) && ({row_reg, col_reg}<16'b0001110111011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001110111011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001110111011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110111011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001110111011011) && ({row_reg, col_reg}<16'b0001110111011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110111011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110111011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110111011111) && ({row_reg, col_reg}<16'b0001110111100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110111100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001110111100011) && ({row_reg, col_reg}<16'b0001110111100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110111100101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001110111100110) && ({row_reg, col_reg}<16'b0001110111101011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110111101011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001110111101100) && ({row_reg, col_reg}<16'b0001110111101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001110111101111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001110111110000) && ({row_reg, col_reg}<16'b0001110111110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001110111110011) && ({row_reg, col_reg}<16'b0001110111110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001110111110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110111110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001110111110111) && ({row_reg, col_reg}<16'b0001110111111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001110111111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001110111111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001110111111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001110111111100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001110111111101)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}>=16'b0001110111111110) && ({row_reg, col_reg}<16'b0001111000000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001111000000000) && ({row_reg, col_reg}<16'b0001111000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111000000101) && ({row_reg, col_reg}<16'b0001111000000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111000000111) && ({row_reg, col_reg}<16'b0001111000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111000001100) && ({row_reg, col_reg}<16'b0001111000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111000010000) && ({row_reg, col_reg}<16'b0001111000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111000010010) && ({row_reg, col_reg}<16'b0001111000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001111000011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111000011010) && ({row_reg, col_reg}<16'b0001111000100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111000100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111000100100) && ({row_reg, col_reg}<16'b0001111000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001111000101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111000101011) && ({row_reg, col_reg}<16'b0001111000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111000110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111000110110) && ({row_reg, col_reg}<16'b0001111000111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001111000111111) && ({row_reg, col_reg}<16'b0001111001000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111001000001) && ({row_reg, col_reg}<16'b0001111001001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111001001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111001001100) && ({row_reg, col_reg}<16'b0001111001010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001111001010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111001010100) && ({row_reg, col_reg}<16'b0001111001011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111001011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111001011110) && ({row_reg, col_reg}<16'b0001111001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001111001100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111001100010) && ({row_reg, col_reg}<16'b0001111001100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111001100101) && ({row_reg, col_reg}<16'b0001111001101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001111001101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111001101001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001111001101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111001101011) && ({row_reg, col_reg}<16'b0001111001101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111001101110) && ({row_reg, col_reg}<16'b0001111001110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001111001110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111001110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001111001110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111001110100) && ({row_reg, col_reg}<16'b0001111001110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001111001110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111001110111) && ({row_reg, col_reg}<16'b0001111001111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001111001111001) && ({row_reg, col_reg}<16'b0001111001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111001111011) && ({row_reg, col_reg}<16'b0001111001111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111001111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111001111111) && ({row_reg, col_reg}<16'b0001111010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111010000010) && ({row_reg, col_reg}<16'b0001111010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001111010010100) && ({row_reg, col_reg}<16'b0001111010011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111010011000) && ({row_reg, col_reg}<16'b0001111010011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111010011010) && ({row_reg, col_reg}<16'b0001111010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111010011111) && ({row_reg, col_reg}<16'b0001111010100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001111010100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111010100011) && ({row_reg, col_reg}<16'b0001111010100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111010100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001111010100110) && ({row_reg, col_reg}<16'b0001111010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111010101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111010101001) && ({row_reg, col_reg}<16'b0001111010101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111010101110) && ({row_reg, col_reg}<16'b0001111010110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111010110011) && ({row_reg, col_reg}<16'b0001111010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111010110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111010110110) && ({row_reg, col_reg}<16'b0001111010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111010111000) && ({row_reg, col_reg}<16'b0001111010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001111010111010) && ({row_reg, col_reg}<16'b0001111010111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111010111101) && ({row_reg, col_reg}<16'b0001111011000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111011000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111011000010) && ({row_reg, col_reg}<16'b0001111011000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001111011000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001111011000101) && ({row_reg, col_reg}<16'b0001111011000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111011000111) && ({row_reg, col_reg}<16'b0001111011001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001111011001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111011001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001111011001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111011001101) && ({row_reg, col_reg}<16'b0001111011001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001111011001111) && ({row_reg, col_reg}<16'b0001111011010001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001111011010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111011010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001111011010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111011010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111011010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001111011010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111011010111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0001111011011000) && ({row_reg, col_reg}<16'b0001111011011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111011011010) && ({row_reg, col_reg}<16'b0001111011011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111011011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111011011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111011011111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111011100000) && ({row_reg, col_reg}<16'b0001111011100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111011100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111011100011) && ({row_reg, col_reg}<16'b0001111011100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111011100101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0001111011100110) && ({row_reg, col_reg}<16'b0001111011101010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111011101010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0001111011101011) && ({row_reg, col_reg}<16'b0001111011101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001111011101111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0001111011110000) && ({row_reg, col_reg}<16'b0001111011110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001111011110011) && ({row_reg, col_reg}<16'b0001111011110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001111011110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111011110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001111011110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111011111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111011111001) && ({row_reg, col_reg}<16'b0001111011111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111011111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111011111100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001111011111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111011111110)) color_data = 12'b001100110010;

		if(({row_reg, col_reg}==16'b0001111011111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0001111100000000) && ({row_reg, col_reg}<16'b0001111100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111100000110) && ({row_reg, col_reg}<16'b0001111100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001111100001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111100001101) && ({row_reg, col_reg}<16'b0001111100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111100010000) && ({row_reg, col_reg}<16'b0001111100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111100010010) && ({row_reg, col_reg}<16'b0001111100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001111100011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111100011010) && ({row_reg, col_reg}<16'b0001111100100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111100100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111100100100) && ({row_reg, col_reg}<16'b0001111100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001111100101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111100101011) && ({row_reg, col_reg}<16'b0001111100110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111100110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111100110111) && ({row_reg, col_reg}<16'b0001111100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001111100111101) && ({row_reg, col_reg}<16'b0001111101000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111101000001) && ({row_reg, col_reg}<16'b0001111101001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111101001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111101001100) && ({row_reg, col_reg}<16'b0001111101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001111101010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111101010100) && ({row_reg, col_reg}<16'b0001111101011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111101011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111101011110) && ({row_reg, col_reg}<16'b0001111101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0001111101100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111101100010) && ({row_reg, col_reg}<16'b0001111101100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111101100101) && ({row_reg, col_reg}<16'b0001111101100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111101100111) && ({row_reg, col_reg}<16'b0001111101101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001111101101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111101101011) && ({row_reg, col_reg}<16'b0001111101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111101101110) && ({row_reg, col_reg}<16'b0001111101110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111101110000) && ({row_reg, col_reg}<16'b0001111101110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111101110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001111101110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111101110100) && ({row_reg, col_reg}<16'b0001111101110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111101110111) && ({row_reg, col_reg}<16'b0001111101111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0001111101111001) && ({row_reg, col_reg}<16'b0001111101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111101111011) && ({row_reg, col_reg}<16'b0001111101111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111101111101) && ({row_reg, col_reg}<16'b0001111110000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001111110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111110000010) && ({row_reg, col_reg}<16'b0001111110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001111110010100) && ({row_reg, col_reg}<16'b0001111110011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111110011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001111110011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111110011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111110011100) && ({row_reg, col_reg}<16'b0001111110011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111110011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111110011111) && ({row_reg, col_reg}<16'b0001111110100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001111110100001) && ({row_reg, col_reg}<16'b0001111110100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0001111110100011) && ({row_reg, col_reg}<16'b0001111110100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111110100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001111110100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001111110100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001111110101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0001111110101001) && ({row_reg, col_reg}<16'b0001111110101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0001111110101110) && ({row_reg, col_reg}<16'b0001111110110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001111110110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001111110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111110110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001111110110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111110110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0001111110111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0001111110111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111110111010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0001111110111011) && ({row_reg, col_reg}<16'b0001111110111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0001111110111110) && ({row_reg, col_reg}<16'b0001111111000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001111111000000) && ({row_reg, col_reg}<16'b0001111111000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111111000010) && ({row_reg, col_reg}<16'b0001111111000100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0001111111000100) && ({row_reg, col_reg}<16'b0001111111000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111111000111) && ({row_reg, col_reg}<16'b0001111111001001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001111111001001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0001111111001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111111001011) && ({row_reg, col_reg}<16'b0001111111001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001111111001101) && ({row_reg, col_reg}<16'b0001111111001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111111001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111111010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0001111111010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0001111111010010) && ({row_reg, col_reg}<16'b0001111111010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111111010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111111010101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0001111111010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001111111010111) && ({row_reg, col_reg}<16'b0001111111011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111111011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001111111011010) && ({row_reg, col_reg}<16'b0001111111011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001111111011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111111011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001111111011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111111011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001111111100000) && ({row_reg, col_reg}<16'b0001111111100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0001111111100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001111111100011) && ({row_reg, col_reg}<16'b0001111111100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111111100101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0001111111100110) && ({row_reg, col_reg}<16'b0001111111101010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111111101010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0001111111101011) && ({row_reg, col_reg}<16'b0001111111101110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0001111111101110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0001111111101111)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0001111111110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0001111111110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0001111111110010) && ({row_reg, col_reg}<16'b0001111111110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0001111111110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111111110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0001111111110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0001111111111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0001111111111001) && ({row_reg, col_reg}<16'b0001111111111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0001111111111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111111111100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0001111111111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0001111111111110)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}==16'b0001111111111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010000000000000) && ({row_reg, col_reg}<16'b0010000000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000000000101) && ({row_reg, col_reg}<16'b0010000000001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010000000001010) && ({row_reg, col_reg}<16'b0010000000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000000001100) && ({row_reg, col_reg}<16'b0010000000001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010000000001110) && ({row_reg, col_reg}<16'b0010000000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000000010000) && ({row_reg, col_reg}<16'b0010000000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000000010010) && ({row_reg, col_reg}<16'b0010000000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010000000011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000000011010) && ({row_reg, col_reg}<16'b0010000000100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000000100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000000100100) && ({row_reg, col_reg}<16'b0010000000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010000000101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000000101011) && ({row_reg, col_reg}<16'b0010000000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000000110100) && ({row_reg, col_reg}<16'b0010000000110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000000110110) && ({row_reg, col_reg}<16'b0010000000111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010000000111110) && ({row_reg, col_reg}<16'b0010000001000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010000001000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000001000010) && ({row_reg, col_reg}<16'b0010000001000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010000001000100) && ({row_reg, col_reg}<16'b0010000001001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000001001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000001001100) && ({row_reg, col_reg}<16'b0010000001010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010000001010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000001010100) && ({row_reg, col_reg}<16'b0010000001011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000001011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000001011110) && ({row_reg, col_reg}<16'b0010000001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010000001100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000001100010) && ({row_reg, col_reg}<16'b0010000001100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000001100101) && ({row_reg, col_reg}<16'b0010000001101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010000001101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000001101001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010000001101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000001101011) && ({row_reg, col_reg}<16'b0010000001101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000001101110) && ({row_reg, col_reg}<16'b0010000001110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000001110000) && ({row_reg, col_reg}<16'b0010000001110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000001110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010000001110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000001110100) && ({row_reg, col_reg}<16'b0010000001110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000001110111) && ({row_reg, col_reg}<16'b0010000001111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010000001111001) && ({row_reg, col_reg}<16'b0010000001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010000001111011) && ({row_reg, col_reg}<16'b0010000001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000001111101) && ({row_reg, col_reg}<16'b0010000010000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000010000010) && ({row_reg, col_reg}<16'b0010000010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010000010010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010000010010101) && ({row_reg, col_reg}<16'b0010000010011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000010011011) && ({row_reg, col_reg}<16'b0010000010011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010000010011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000010011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010000010011111) && ({row_reg, col_reg}<16'b0010000010100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010000010100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000010100010) && ({row_reg, col_reg}<16'b0010000010100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000010100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010000010100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010000010100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010000010101000) && ({row_reg, col_reg}<16'b0010000010101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000010101011) && ({row_reg, col_reg}<16'b0010000010101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010000010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000010101110) && ({row_reg, col_reg}<16'b0010000010110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000010110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000010110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000010110110) && ({row_reg, col_reg}<16'b0010000010111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000010111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010000010111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010000010111011) && ({row_reg, col_reg}<16'b0010000010111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010000010111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010000010111110) && ({row_reg, col_reg}<16'b0010000011000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000011000001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010000011000010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010000011000011) && ({row_reg, col_reg}<16'b0010000011000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000011000111) && ({row_reg, col_reg}<16'b0010000011001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010000011001001) && ({row_reg, col_reg}<16'b0010000011001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000011001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000011001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000011001101) && ({row_reg, col_reg}<16'b0010000011010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000011010000) && ({row_reg, col_reg}<16'b0010000011010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010000011010010) && ({row_reg, col_reg}<16'b0010000011010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000011010101) && ({row_reg, col_reg}<16'b0010000011010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000011010111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010000011011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000011011001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010000011011010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010000011011011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010000011011100) && ({row_reg, col_reg}<16'b0010000011011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000011011110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010000011011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000011100000) && ({row_reg, col_reg}<16'b0010000011100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000011100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000011100100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010000011100101) && ({row_reg, col_reg}<16'b0010000011101010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000011101010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010000011101011) && ({row_reg, col_reg}<16'b0010000011101110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010000011101110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0010000011101111) && ({row_reg, col_reg}<16'b0010000011110001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010000011110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000011110010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010000011110011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010000011110100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010000011110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000011110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000011110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010000011111000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0010000011111001) && ({row_reg, col_reg}<16'b0010000011111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000011111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000011111100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010000011111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000011111110)) color_data = 12'b001100110001;

		if(({row_reg, col_reg}==16'b0010000011111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000100000000) && ({row_reg, col_reg}<16'b0010000100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000100000101) && ({row_reg, col_reg}<16'b0010000100001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000100001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010000100001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000100001010) && ({row_reg, col_reg}<16'b0010000100001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000100001100) && ({row_reg, col_reg}<16'b0010000100001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010000100001110) && ({row_reg, col_reg}<16'b0010000100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000100010010) && ({row_reg, col_reg}<16'b0010000100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010000100011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000100011010) && ({row_reg, col_reg}<16'b0010000100100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000100100010) && ({row_reg, col_reg}<16'b0010000100100100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000100100100) && ({row_reg, col_reg}<16'b0010000100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010000100101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000100101011) && ({row_reg, col_reg}<16'b0010000100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000100110100) && ({row_reg, col_reg}<16'b0010000100110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000100110110) && ({row_reg, col_reg}<16'b0010000100111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010000100111110) && ({row_reg, col_reg}<16'b0010000101000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000101000001) && ({row_reg, col_reg}<16'b0010000101000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010000101000100) && ({row_reg, col_reg}<16'b0010000101001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000101001010) && ({row_reg, col_reg}<16'b0010000101001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000101001100) && ({row_reg, col_reg}<16'b0010000101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010000101010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000101010100) && ({row_reg, col_reg}<16'b0010000101011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000101011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000101011110) && ({row_reg, col_reg}<16'b0010000101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010000101100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000101100010) && ({row_reg, col_reg}<16'b0010000101100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000101100101) && ({row_reg, col_reg}<16'b0010000101101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000101101000) && ({row_reg, col_reg}<16'b0010000101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000101101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000101101011) && ({row_reg, col_reg}<16'b0010000101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000101101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000101101111) && ({row_reg, col_reg}<16'b0010000101110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000101110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000101110011) && ({row_reg, col_reg}<16'b0010000101110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000101110111) && ({row_reg, col_reg}<16'b0010000101111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010000101111001) && ({row_reg, col_reg}<16'b0010000101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010000101111011) && ({row_reg, col_reg}<16'b0010000101111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000101111101) && ({row_reg, col_reg}<16'b0010000110000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000110000010) && ({row_reg, col_reg}<16'b0010000110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010000110010100) && ({row_reg, col_reg}<16'b0010000110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000110010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000110011000) && ({row_reg, col_reg}<16'b0010000110011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010000110011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000110011011) && ({row_reg, col_reg}<16'b0010000110011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010000110011101) && ({row_reg, col_reg}<16'b0010000110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000110011111) && ({row_reg, col_reg}<16'b0010000110100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010000110100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010000110100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000110100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010000110100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000110100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010000110100110) && ({row_reg, col_reg}<16'b0010000110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010000110101000) && ({row_reg, col_reg}<16'b0010000110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000110101010) && ({row_reg, col_reg}<16'b0010000110101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010000110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010000110101110) && ({row_reg, col_reg}<16'b0010000110110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010000110110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010000110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000110110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010000110110110) && ({row_reg, col_reg}<16'b0010000110111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010000110111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010000110111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010000110111010) && ({row_reg, col_reg}<16'b0010000110111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010000110111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010000110111101) && ({row_reg, col_reg}<16'b0010000111000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000111000001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010000111000010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010000111000011) && ({row_reg, col_reg}<16'b0010000111000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000111000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010000111000110) && ({row_reg, col_reg}<16'b0010000111001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000111001000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010000111001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000111001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010000111001011) && ({row_reg, col_reg}<16'b0010000111001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010000111001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000111001110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010000111001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010000111010000) && ({row_reg, col_reg}<16'b0010000111010010)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0010000111010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010000111010011) && ({row_reg, col_reg}<16'b0010000111010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000111010101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010000111010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000111010111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010000111011000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010000111011001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010000111011010)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0010000111011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010000111011100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010000111011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000111011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010000111011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000111100000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010000111100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010000111100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010000111100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000111100100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0010000111100101) && ({row_reg, col_reg}<16'b0010000111101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010000111101110) && ({row_reg, col_reg}<16'b0010000111110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010000111110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010000111110001) && ({row_reg, col_reg}<16'b0010000111110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000111110011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010000111110100) && ({row_reg, col_reg}<16'b0010000111110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000111110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000111110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010000111111000) && ({row_reg, col_reg}<16'b0010000111111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010000111111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010000111111100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010000111111101)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}>=16'b0010000111111110) && ({row_reg, col_reg}<16'b0010001000000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010001000000000) && ({row_reg, col_reg}<16'b0010001000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001000000101) && ({row_reg, col_reg}<16'b0010001000000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010001000000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010001000001000) && ({row_reg, col_reg}<16'b0010001000001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010001000001010) && ({row_reg, col_reg}<16'b0010001000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001000001101) && ({row_reg, col_reg}<16'b0010001000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001000010010) && ({row_reg, col_reg}<16'b0010001000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010001000011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001000011010) && ({row_reg, col_reg}<16'b0010001000100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001000100001) && ({row_reg, col_reg}<16'b0010001000100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001000100011) && ({row_reg, col_reg}<16'b0010001000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010001000101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001000101011) && ({row_reg, col_reg}<16'b0010001000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001000110100) && ({row_reg, col_reg}<16'b0010001000110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001000110110) && ({row_reg, col_reg}<16'b0010001000111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010001000111101) && ({row_reg, col_reg}<16'b0010001001000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001001000001) && ({row_reg, col_reg}<16'b0010001001001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001001001010) && ({row_reg, col_reg}<16'b0010001001001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001001001100) && ({row_reg, col_reg}<16'b0010001001010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010001001010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001001010100) && ({row_reg, col_reg}<16'b0010001001011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001001011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001001011110) && ({row_reg, col_reg}<16'b0010001001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010001001100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001001100010) && ({row_reg, col_reg}<16'b0010001001100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001001100100) && ({row_reg, col_reg}<16'b0010001001101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001001101000) && ({row_reg, col_reg}<16'b0010001001101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001001101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001001101011) && ({row_reg, col_reg}<16'b0010001001101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001001101101) && ({row_reg, col_reg}<16'b0010001001101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001001101111) && ({row_reg, col_reg}<16'b0010001001110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001001110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001001110011) && ({row_reg, col_reg}<16'b0010001001110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001001110111) && ({row_reg, col_reg}<16'b0010001001111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010001001111001) && ({row_reg, col_reg}<16'b0010001001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001001111011) && ({row_reg, col_reg}<16'b0010001001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001001111101) && ({row_reg, col_reg}<16'b0010001010000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010001010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001010000010) && ({row_reg, col_reg}<16'b0010001010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010001010010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001010010101) && ({row_reg, col_reg}<16'b0010001010010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001010010111) && ({row_reg, col_reg}<16'b0010001010011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001010011101) && ({row_reg, col_reg}<16'b0010001010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001010011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010001010100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010001010100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010001010100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001010100011) && ({row_reg, col_reg}<16'b0010001010100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010001010100101) && ({row_reg, col_reg}<16'b0010001010100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001010100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001010101000) && ({row_reg, col_reg}<16'b0010001010101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001010101011) && ({row_reg, col_reg}<16'b0010001010101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010001010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001010101110) && ({row_reg, col_reg}<16'b0010001010110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001010110011) && ({row_reg, col_reg}<16'b0010001010110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001010110110) && ({row_reg, col_reg}<16'b0010001010111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001010111000) && ({row_reg, col_reg}<16'b0010001010111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001010111010) && ({row_reg, col_reg}<16'b0010001010111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001010111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001010111101) && ({row_reg, col_reg}<16'b0010001011000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001011000001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010001011000010) && ({row_reg, col_reg}<16'b0010001011000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001011000101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010001011000110) && ({row_reg, col_reg}<16'b0010001011001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001011001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001011001010) && ({row_reg, col_reg}<16'b0010001011001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010001011001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010001011001110) && ({row_reg, col_reg}<16'b0010001011010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010001011010000) && ({row_reg, col_reg}<16'b0010001011010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010001011010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001011010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010001011010100) && ({row_reg, col_reg}<16'b0010001011010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001011010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010001011010111) && ({row_reg, col_reg}<16'b0010001011011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001011011001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010001011011010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0010001011011011)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0010001011011100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010001011011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001011011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010001011011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001011100000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001011100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010001011100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001011100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010001011100100) && ({row_reg, col_reg}<16'b0010001011100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010001011100111) && ({row_reg, col_reg}<16'b0010001011101001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010001011101001) && ({row_reg, col_reg}<16'b0010001011101011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010001011101011) && ({row_reg, col_reg}<16'b0010001011101110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001011101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010001011101111) && ({row_reg, col_reg}<16'b0010001011110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001011110001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010001011110010) && ({row_reg, col_reg}<16'b0010001011110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010001011110110) && ({row_reg, col_reg}<16'b0010001011111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010001011111000) && ({row_reg, col_reg}<16'b0010001011111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001011111101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001011111110)) color_data = 12'b001100100010;

		if(({row_reg, col_reg}==16'b0010001011111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010001100000000) && ({row_reg, col_reg}<16'b0010001100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001100000101) && ({row_reg, col_reg}<16'b0010001100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010001100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010001100001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010001100001010) && ({row_reg, col_reg}<16'b0010001100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001100010010) && ({row_reg, col_reg}<16'b0010001100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010001100011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001100011010) && ({row_reg, col_reg}<16'b0010001100100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001100100001) && ({row_reg, col_reg}<16'b0010001100100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001100100011) && ({row_reg, col_reg}<16'b0010001100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010001100101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001100101011) && ({row_reg, col_reg}<16'b0010001100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001100110100) && ({row_reg, col_reg}<16'b0010001100110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001100110110) && ({row_reg, col_reg}<16'b0010001101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010001101000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001101000001) && ({row_reg, col_reg}<16'b0010001101001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001101001010) && ({row_reg, col_reg}<16'b0010001101001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001101001100) && ({row_reg, col_reg}<16'b0010001101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010001101010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001101010100) && ({row_reg, col_reg}<16'b0010001101011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001101011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001101011110) && ({row_reg, col_reg}<16'b0010001101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010001101100001) && ({row_reg, col_reg}<16'b0010001101100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001101100100) && ({row_reg, col_reg}<16'b0010001101101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001101101000) && ({row_reg, col_reg}<16'b0010001101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001101101010) && ({row_reg, col_reg}<16'b0010001101101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001101101100) && ({row_reg, col_reg}<16'b0010001101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001101101110) && ({row_reg, col_reg}<16'b0010001101110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010001101110000) && ({row_reg, col_reg}<16'b0010001101110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001101110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010001101110011) && ({row_reg, col_reg}<16'b0010001101110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001101110111) && ({row_reg, col_reg}<16'b0010001101111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010001101111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001101111011) && ({row_reg, col_reg}<16'b0010001101111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001101111101) && ({row_reg, col_reg}<16'b0010001110000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010001110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001110000010) && ({row_reg, col_reg}<16'b0010001110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010001110010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001110010101) && ({row_reg, col_reg}<16'b0010001110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010001110010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001110011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001110011001) && ({row_reg, col_reg}<16'b0010001110011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001110011101) && ({row_reg, col_reg}<16'b0010001110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001110011111) && ({row_reg, col_reg}<16'b0010001110100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010001110100001) && ({row_reg, col_reg}<16'b0010001110100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010001110100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001110100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010001110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001110100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001110101000) && ({row_reg, col_reg}<16'b0010001110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010001110101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010001110101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010001110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001110101110) && ({row_reg, col_reg}<16'b0010001110110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010001110110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010001110110011) && ({row_reg, col_reg}<16'b0010001110110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010001110110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010001110110110) && ({row_reg, col_reg}<16'b0010001110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010001110111000) && ({row_reg, col_reg}<16'b0010001110111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010001110111011) && ({row_reg, col_reg}<16'b0010001110111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010001110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001110111110) && ({row_reg, col_reg}<16'b0010001111000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001111000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010001111000010) && ({row_reg, col_reg}<16'b0010001111000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010001111000100) && ({row_reg, col_reg}<16'b0010001111000110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001111000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010001111000111) && ({row_reg, col_reg}<16'b0010001111001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001111001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010001111001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010001111001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010001111001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010001111001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001111001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001111001111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010001111010000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0010001111010001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0010001111010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010001111010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010001111010100) && ({row_reg, col_reg}<16'b0010001111010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001111010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001111010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010001111011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001111011001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0010001111011010) && ({row_reg, col_reg}<16'b0010001111011101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010001111011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001111011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010001111011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010001111100000) && ({row_reg, col_reg}<16'b0010001111100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010001111100010) && ({row_reg, col_reg}<16'b0010001111100100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010001111100100) && ({row_reg, col_reg}<16'b0010001111100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001111100110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010001111100111) && ({row_reg, col_reg}<16'b0010001111101001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010001111101001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010001111101010) && ({row_reg, col_reg}<16'b0010001111101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001111101100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010001111101101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0010001111101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001111101111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010001111110000) && ({row_reg, col_reg}<16'b0010001111110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010001111110010) && ({row_reg, col_reg}<16'b0010001111110100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001111110100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010001111110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001111110110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010001111110111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010001111111000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010001111111001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010001111111010) && ({row_reg, col_reg}<16'b0010001111111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010001111111101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010001111111110)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}==16'b0010001111111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010000000000) && ({row_reg, col_reg}<16'b0010010000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010000000101) && ({row_reg, col_reg}<16'b0010010000000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010000000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010010000001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010010000001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010000001011) && ({row_reg, col_reg}<16'b0010010000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010000010010) && ({row_reg, col_reg}<16'b0010010000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010010000011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010000011010) && ({row_reg, col_reg}<16'b0010010000100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010000100001) && ({row_reg, col_reg}<16'b0010010000100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010000100011) && ({row_reg, col_reg}<16'b0010010000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010010000101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010000101011) && ({row_reg, col_reg}<16'b0010010000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010000110100) && ({row_reg, col_reg}<16'b0010010000110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010000110110) && ({row_reg, col_reg}<16'b0010010001000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010010001000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010001000001) && ({row_reg, col_reg}<16'b0010010001001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010001001010) && ({row_reg, col_reg}<16'b0010010001001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010001001100) && ({row_reg, col_reg}<16'b0010010001010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010010001010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010001010100) && ({row_reg, col_reg}<16'b0010010001011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010001011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010001011110) && ({row_reg, col_reg}<16'b0010010001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010010001100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010001100010) && ({row_reg, col_reg}<16'b0010010001100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010010001100101) && ({row_reg, col_reg}<16'b0010010001101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010001101000) && ({row_reg, col_reg}<16'b0010010001101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010001101010) && ({row_reg, col_reg}<16'b0010010001101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010001101101) && ({row_reg, col_reg}<16'b0010010001101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010001101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010010001110000) && ({row_reg, col_reg}<16'b0010010001110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010001110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010001110011) && ({row_reg, col_reg}<16'b0010010001110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010001110111) && ({row_reg, col_reg}<16'b0010010001111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010010001111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010001111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010010001111011) && ({row_reg, col_reg}<16'b0010010001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010001111101) && ({row_reg, col_reg}<16'b0010010010000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010010000010) && ({row_reg, col_reg}<16'b0010010010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010010010010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010010010101) && ({row_reg, col_reg}<16'b0010010010011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010010011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010010011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010010010011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010010010011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010010011101) && ({row_reg, col_reg}<16'b0010010010100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010010100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010010100001) && ({row_reg, col_reg}<16'b0010010010100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010010100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010010010100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010010010100101) && ({row_reg, col_reg}<16'b0010010010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010010101000) && ({row_reg, col_reg}<16'b0010010010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010010101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010010010101011) && ({row_reg, col_reg}<16'b0010010010101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010010101101) && ({row_reg, col_reg}<16'b0010010010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010010010110010) && ({row_reg, col_reg}<16'b0010010010110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010010010110100) && ({row_reg, col_reg}<16'b0010010010110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010010110110) && ({row_reg, col_reg}<16'b0010010010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010010111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010010111011) && ({row_reg, col_reg}<16'b0010010010111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010010010111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010010111110) && ({row_reg, col_reg}<16'b0010010011000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010011000001) && ({row_reg, col_reg}<16'b0010010011000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010011000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010011000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010011000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010011000111) && ({row_reg, col_reg}<16'b0010010011001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010011001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010011001110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010010011001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010011010000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0010010011010001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010010011010010)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0010010011010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010010011010100) && ({row_reg, col_reg}<16'b0010010011010110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010010011010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010011010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010011011000)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0010010011011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010010011011010) && ({row_reg, col_reg}<16'b0010010011011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010011011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010010011011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010011011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010010011011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010011100000) && ({row_reg, col_reg}<16'b0010010011100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010011100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010011100011) && ({row_reg, col_reg}<16'b0010010011100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010011100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010010011100110) && ({row_reg, col_reg}<16'b0010010011101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010010011101010) && ({row_reg, col_reg}<16'b0010010011101100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010010011101100) && ({row_reg, col_reg}<16'b0010010011101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010010011101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010010011110000) && ({row_reg, col_reg}<16'b0010010011110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010011110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010011110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010011110100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010010011110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010010011110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010011110111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0010010011111000) && ({row_reg, col_reg}<16'b0010010011111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010010011111010) && ({row_reg, col_reg}<16'b0010010011111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010011111101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010011111110)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}==16'b0010010011111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010100000000) && ({row_reg, col_reg}<16'b0010010100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010100000101) && ({row_reg, col_reg}<16'b0010010100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010010100001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010010100001010) && ({row_reg, col_reg}<16'b0010010100001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010100001100) && ({row_reg, col_reg}<16'b0010010100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010100010000) && ({row_reg, col_reg}<16'b0010010100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010100010010) && ({row_reg, col_reg}<16'b0010010100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010010100011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010100011010) && ({row_reg, col_reg}<16'b0010010100100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010100100011) && ({row_reg, col_reg}<16'b0010010100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010010100101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010100101011) && ({row_reg, col_reg}<16'b0010010100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010100110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010100110110) && ({row_reg, col_reg}<16'b0010010101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010010101000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010101000001) && ({row_reg, col_reg}<16'b0010010101000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010010101000101) && ({row_reg, col_reg}<16'b0010010101001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010101001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010101001100) && ({row_reg, col_reg}<16'b0010010101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010010101010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010101010100) && ({row_reg, col_reg}<16'b0010010101011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010101011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010101011110) && ({row_reg, col_reg}<16'b0010010101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010010101100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010101100010) && ({row_reg, col_reg}<16'b0010010101100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010010101100101) && ({row_reg, col_reg}<16'b0010010101101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010101101000) && ({row_reg, col_reg}<16'b0010010101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010101101010) && ({row_reg, col_reg}<16'b0010010101101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010101101101) && ({row_reg, col_reg}<16'b0010010101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010101101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010010101110000) && ({row_reg, col_reg}<16'b0010010101110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010101110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010101110011) && ({row_reg, col_reg}<16'b0010010101110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010101110111) && ({row_reg, col_reg}<16'b0010010101111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010010101111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010101111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010101111011) && ({row_reg, col_reg}<16'b0010010101111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010101111101) && ({row_reg, col_reg}<16'b0010010110000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010110000010) && ({row_reg, col_reg}<16'b0010010110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010010110010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010110010101) && ({row_reg, col_reg}<16'b0010010110011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010110011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010010110011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010110011011) && ({row_reg, col_reg}<16'b0010010110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010010110011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010010110011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010010110011111) && ({row_reg, col_reg}<16'b0010010110100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010010110100001) && ({row_reg, col_reg}<16'b0010010110100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010010110100011) && ({row_reg, col_reg}<16'b0010010110100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010010110100101) && ({row_reg, col_reg}<16'b0010010110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010110101000) && ({row_reg, col_reg}<16'b0010010110101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010010110101011) && ({row_reg, col_reg}<16'b0010010110101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010110101101) && ({row_reg, col_reg}<16'b0010010110110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010110110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010010110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010110110100) && ({row_reg, col_reg}<16'b0010010110110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010010110110110) && ({row_reg, col_reg}<16'b0010010110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010010110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010110111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010110111011) && ({row_reg, col_reg}<16'b0010010110111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010010110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010010110111110) && ({row_reg, col_reg}<16'b0010010111000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010111000001) && ({row_reg, col_reg}<16'b0010010111000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010111000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010010111000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010010111000110) && ({row_reg, col_reg}<16'b0010010111001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010111001000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010010111001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010010111001010) && ({row_reg, col_reg}<16'b0010010111001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010111001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010111001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010010111010000) && ({row_reg, col_reg}<16'b0010010111010011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010010111010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010111010100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010010111010101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010010111010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010111010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010111011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010010111011001)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0010010111011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010010111011011) && ({row_reg, col_reg}<16'b0010010111011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010111011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010010111011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010111100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010010111100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010111100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010010111100011) && ({row_reg, col_reg}<16'b0010010111100110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010010111100110) && ({row_reg, col_reg}<16'b0010010111101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010010111101010) && ({row_reg, col_reg}<16'b0010010111101100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010010111101100) && ({row_reg, col_reg}<16'b0010010111101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010010111101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010111110000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010010111110001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010010111110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010010111110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010111110100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010010111110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010010111110110) && ({row_reg, col_reg}<16'b0010010111111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010010111111000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010010111111001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010010111111010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010010111111011) && ({row_reg, col_reg}<16'b0010010111111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010010111111110)) color_data = 12'b001100100010;

		if(({row_reg, col_reg}==16'b0010010111111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011000000000) && ({row_reg, col_reg}<16'b0010011000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011000000101) && ({row_reg, col_reg}<16'b0010011000000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010011000000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010011000001000) && ({row_reg, col_reg}<16'b0010011000001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010011000001010) && ({row_reg, col_reg}<16'b0010011000001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011000001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010011000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011000010000) && ({row_reg, col_reg}<16'b0010011000010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011000010010) && ({row_reg, col_reg}<16'b0010011000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011000011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011000011010) && ({row_reg, col_reg}<16'b0010011000100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011000100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011000100100) && ({row_reg, col_reg}<16'b0010011000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011000101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011000101011) && ({row_reg, col_reg}<16'b0010011000110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011000110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011000110111) && ({row_reg, col_reg}<16'b0010011000111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010011000111101) && ({row_reg, col_reg}<16'b0010011001000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011001000001) && ({row_reg, col_reg}<16'b0010011001000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011001000100) && ({row_reg, col_reg}<16'b0010011001000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010011001000110) && ({row_reg, col_reg}<16'b0010011001001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011001001100) && ({row_reg, col_reg}<16'b0010011001010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011001010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011001010100) && ({row_reg, col_reg}<16'b0010011001011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011001011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011001011110) && ({row_reg, col_reg}<16'b0010011001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011001100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011001100010) && ({row_reg, col_reg}<16'b0010011001100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010011001100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011001100101) && ({row_reg, col_reg}<16'b0010011001101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010011001101000) && ({row_reg, col_reg}<16'b0010011001101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011001101010) && ({row_reg, col_reg}<16'b0010011001101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010011001101100) && ({row_reg, col_reg}<16'b0010011001101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011001101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010011001101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010011001110000) && ({row_reg, col_reg}<16'b0010011001110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011001110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011001110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011001110100) && ({row_reg, col_reg}<16'b0010011001110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011001110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010011001111000) && ({row_reg, col_reg}<16'b0010011001111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011001111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010011001111011) && ({row_reg, col_reg}<16'b0010011001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011001111101) && ({row_reg, col_reg}<16'b0010011010000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010011010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011010000010) && ({row_reg, col_reg}<16'b0010011010010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010011010010101) && ({row_reg, col_reg}<16'b0010011010011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010011010011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011010011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011010011011) && ({row_reg, col_reg}<16'b0010011010011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011010011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010011010011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011010011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011010100000) && ({row_reg, col_reg}<16'b0010011010100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010011010100010) && ({row_reg, col_reg}<16'b0010011010100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010011010100101) && ({row_reg, col_reg}<16'b0010011010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011010101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010011010101001) && ({row_reg, col_reg}<16'b0010011010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011010101101) && ({row_reg, col_reg}<16'b0010011010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010011010110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010011010110011) && ({row_reg, col_reg}<16'b0010011010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011010110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011010110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010011010111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010011010111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011010111010) && ({row_reg, col_reg}<16'b0010011010111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011010111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010011010111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011010111110) && ({row_reg, col_reg}<16'b0010011011000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010011011000001) && ({row_reg, col_reg}<16'b0010011011000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011011000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011011000101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010011011000110) && ({row_reg, col_reg}<16'b0010011011001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010011011001000) && ({row_reg, col_reg}<16'b0010011011001010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011011001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010011011001011) && ({row_reg, col_reg}<16'b0010011011001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011011001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011011001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010011011010000) && ({row_reg, col_reg}<16'b0010011011010011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010011011010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011011010100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010011011010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011011010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011011010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010011011011000) && ({row_reg, col_reg}<16'b0010011011011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011011011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010011011011011) && ({row_reg, col_reg}<16'b0010011011011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010011011011110) && ({row_reg, col_reg}<16'b0010011011100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011011100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011011100010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010011011100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010011011100100) && ({row_reg, col_reg}<16'b0010011011100110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010011011100110) && ({row_reg, col_reg}<16'b0010011011101000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010011011101000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0010011011101001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010011011101010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010011011101011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010011011101100) && ({row_reg, col_reg}<16'b0010011011101110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010011011101110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010011011101111) && ({row_reg, col_reg}<16'b0010011011110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011011110001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010011011110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010011011110011) && ({row_reg, col_reg}<16'b0010011011110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010011011110110) && ({row_reg, col_reg}<16'b0010011011111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011011111000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011011111001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010011011111010) && ({row_reg, col_reg}<16'b0010011011111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011011111110)) color_data = 12'b001100100010;

		if(({row_reg, col_reg}==16'b0010011011111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011100000000) && ({row_reg, col_reg}<16'b0010011100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011100000101) && ({row_reg, col_reg}<16'b0010011100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010011100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010011100001000) && ({row_reg, col_reg}<16'b0010011100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010011100001010) && ({row_reg, col_reg}<16'b0010011100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011100010010) && ({row_reg, col_reg}<16'b0010011100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011100011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011100011010) && ({row_reg, col_reg}<16'b0010011100100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011100100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010011100100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011100100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011100100100) && ({row_reg, col_reg}<16'b0010011100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011100101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011100101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010011100101100) && ({row_reg, col_reg}<16'b0010011100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010011100110001) && ({row_reg, col_reg}<16'b0010011100110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011100110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011100110111) && ({row_reg, col_reg}<16'b0010011100111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010011100111110) && ({row_reg, col_reg}<16'b0010011101000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011101000001) && ({row_reg, col_reg}<16'b0010011101000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010011101000100) && ({row_reg, col_reg}<16'b0010011101001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011101001001) && ({row_reg, col_reg}<16'b0010011101001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010011101001100) && ({row_reg, col_reg}<16'b0010011101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011101010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011101010100) && ({row_reg, col_reg}<16'b0010011101011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011101011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011101011110) && ({row_reg, col_reg}<16'b0010011101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010011101100001) && ({row_reg, col_reg}<16'b0010011101100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011101100100) && ({row_reg, col_reg}<16'b0010011101101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010011101101000) && ({row_reg, col_reg}<16'b0010011101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011101101010) && ({row_reg, col_reg}<16'b0010011101101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010011101101100) && ({row_reg, col_reg}<16'b0010011101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010011101101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010011101110000) && ({row_reg, col_reg}<16'b0010011101110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011101110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011101110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011101110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011101110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011101110110) && ({row_reg, col_reg}<16'b0010011101111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010011101111000) && ({row_reg, col_reg}<16'b0010011101111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011101111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010011101111011) && ({row_reg, col_reg}<16'b0010011101111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011101111101) && ({row_reg, col_reg}<16'b0010011110000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010011110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011110000010) && ({row_reg, col_reg}<16'b0010011110010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010011110010101) && ({row_reg, col_reg}<16'b0010011110010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011110010111) && ({row_reg, col_reg}<16'b0010011110011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010011110011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010011110011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010011110011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010011110011101) && ({row_reg, col_reg}<16'b0010011110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011110011111) && ({row_reg, col_reg}<16'b0010011110100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010011110100010) && ({row_reg, col_reg}<16'b0010011110100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010011110100101) && ({row_reg, col_reg}<16'b0010011110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011110101000) && ({row_reg, col_reg}<16'b0010011110101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010011110101110) && ({row_reg, col_reg}<16'b0010011110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010011110110000) && ({row_reg, col_reg}<16'b0010011110110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010011110110011) && ({row_reg, col_reg}<16'b0010011110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011110110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011110110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010011110110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010011110111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010011110111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011110111010) && ({row_reg, col_reg}<16'b0010011110111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010011110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011110111110) && ({row_reg, col_reg}<16'b0010011111000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010011111000001) && ({row_reg, col_reg}<16'b0010011111000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010011111000100) && ({row_reg, col_reg}<16'b0010011111001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011111001000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011111001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010011111001010) && ({row_reg, col_reg}<16'b0010011111001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011111001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011111001110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010011111001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011111010000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010011111010001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010011111010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010011111010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011111010100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010011111010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011111010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010011111010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010011111011000) && ({row_reg, col_reg}<16'b0010011111011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010011111011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010011111011011) && ({row_reg, col_reg}<16'b0010011111011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011111011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010011111011110) && ({row_reg, col_reg}<16'b0010011111100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011111100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010011111100001) && ({row_reg, col_reg}<16'b0010011111100100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010011111100100) && ({row_reg, col_reg}<16'b0010011111100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011111100111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010011111101000)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}>=16'b0010011111101001) && ({row_reg, col_reg}<16'b0010011111101011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010011111101011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011111101100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010011111101101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010011111101110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010011111101111) && ({row_reg, col_reg}<16'b0010011111110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011111110001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010011111110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011111110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011111110100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010011111110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010011111110110) && ({row_reg, col_reg}<16'b0010011111111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010011111111000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010011111111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011111111010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010011111111011) && ({row_reg, col_reg}<16'b0010011111111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010011111111101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010011111111110)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}==16'b0010011111111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010100000000000) && ({row_reg, col_reg}<16'b0010100000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100000000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010100000000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010100000000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010100000001000) && ({row_reg, col_reg}<16'b0010100000001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100000001101) && ({row_reg, col_reg}<16'b0010100000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100000010010) && ({row_reg, col_reg}<16'b0010100000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100000011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100000011010) && ({row_reg, col_reg}<16'b0010100000100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100000100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010100000100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100000100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100000100100) && ({row_reg, col_reg}<16'b0010100000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010100000101010) && ({row_reg, col_reg}<16'b0010100000101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100000101100) && ({row_reg, col_reg}<16'b0010100000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100000110000) && ({row_reg, col_reg}<16'b0010100000110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100000110010) && ({row_reg, col_reg}<16'b0010100000110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100000110100) && ({row_reg, col_reg}<16'b0010100000110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100000110110) && ({row_reg, col_reg}<16'b0010100000111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010100000111110) && ({row_reg, col_reg}<16'b0010100001000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010100001000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100001000010) && ({row_reg, col_reg}<16'b0010100001000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100001000100) && ({row_reg, col_reg}<16'b0010100001001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100001001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100001001100) && ({row_reg, col_reg}<16'b0010100001010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100001010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100001010100) && ({row_reg, col_reg}<16'b0010100001011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100001011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100001011110) && ({row_reg, col_reg}<16'b0010100001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010100001100001) && ({row_reg, col_reg}<16'b0010100001100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100001100011) && ({row_reg, col_reg}<16'b0010100001100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100001100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010100001101000) && ({row_reg, col_reg}<16'b0010100001101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100001101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010100001101011) && ({row_reg, col_reg}<16'b0010100001101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100001101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010100001101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010100001110000) && ({row_reg, col_reg}<16'b0010100001110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100001110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100001110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100001110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100001110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100001110110) && ({row_reg, col_reg}<16'b0010100001111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010100001111000) && ({row_reg, col_reg}<16'b0010100001111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100001111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010100001111011) && ({row_reg, col_reg}<16'b0010100001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100001111101) && ({row_reg, col_reg}<16'b0010100010000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010100010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100010000010) && ({row_reg, col_reg}<16'b0010100010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100010010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100010010101) && ({row_reg, col_reg}<16'b0010100010011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100010011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010100010011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010100010011100) && ({row_reg, col_reg}<16'b0010100010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100010011111) && ({row_reg, col_reg}<16'b0010100010100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010100010100001) && ({row_reg, col_reg}<16'b0010100010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100010100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100010100101) && ({row_reg, col_reg}<16'b0010100010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010100010101000) && ({row_reg, col_reg}<16'b0010100010101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100010101011) && ({row_reg, col_reg}<16'b0010100010101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100010101110) && ({row_reg, col_reg}<16'b0010100010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100010110000) && ({row_reg, col_reg}<16'b0010100010110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010100010110011) && ({row_reg, col_reg}<16'b0010100010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100010110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100010110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010100010111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010100010111001) && ({row_reg, col_reg}<16'b0010100010111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100010111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010100010111100) && ({row_reg, col_reg}<16'b0010100010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010100010111110) && ({row_reg, col_reg}<16'b0010100011000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010100011000010) && ({row_reg, col_reg}<16'b0010100011000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010100011000100) && ({row_reg, col_reg}<16'b0010100011001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010100011001000) && ({row_reg, col_reg}<16'b0010100011001010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010100011001010) && ({row_reg, col_reg}<16'b0010100011001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010100011001110) && ({row_reg, col_reg}<16'b0010100011010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100011010000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0010100011010001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010100011010010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0010100011010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100011010100) && ({row_reg, col_reg}<16'b0010100011010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100011010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010100011010111) && ({row_reg, col_reg}<16'b0010100011011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100011011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100011011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010100011011011) && ({row_reg, col_reg}<16'b0010100011011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100011011101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010100011011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100011011111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010100011100000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010100011100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010100011100010) && ({row_reg, col_reg}<16'b0010100011100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100011100110)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0010100011100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010100011101000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0010100011101001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010100011101010)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0010100011101011) && ({row_reg, col_reg}<16'b0010100011101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100011101101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010100011101110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010100011101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010100011110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100011110001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010100011110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010100011110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100011110100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010100011110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100011110110) && ({row_reg, col_reg}<16'b0010100011111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100011111000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010100011111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100011111010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010100011111011) && ({row_reg, col_reg}<16'b0010100011111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100011111101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010100011111110)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}==16'b0010100011111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010100100000000) && ({row_reg, col_reg}<16'b0010100100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100100000101) && ({row_reg, col_reg}<16'b0010100100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010100100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010100100001000) && ({row_reg, col_reg}<16'b0010100100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100100001100) && ({row_reg, col_reg}<16'b0010100100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100100010010) && ({row_reg, col_reg}<16'b0010100100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100100011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100100011010) && ({row_reg, col_reg}<16'b0010100100100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100100100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100100100100) && ({row_reg, col_reg}<16'b0010100100101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100100101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100100101010) && ({row_reg, col_reg}<16'b0010100100101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100100101100) && ({row_reg, col_reg}<16'b0010100100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100100110000) && ({row_reg, col_reg}<16'b0010100100110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100100110010) && ({row_reg, col_reg}<16'b0010100100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100100110100) && ({row_reg, col_reg}<16'b0010100100110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100100110110) && ({row_reg, col_reg}<16'b0010100100111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010100100111110) && ({row_reg, col_reg}<16'b0010100101000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010100101000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100101000010) && ({row_reg, col_reg}<16'b0010100101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100101000100) && ({row_reg, col_reg}<16'b0010100101001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100101001010) && ({row_reg, col_reg}<16'b0010100101001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100101001100) && ({row_reg, col_reg}<16'b0010100101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100101010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100101010100) && ({row_reg, col_reg}<16'b0010100101011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100101011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100101011110) && ({row_reg, col_reg}<16'b0010100101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010100101100001) && ({row_reg, col_reg}<16'b0010100101100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100101100100) && ({row_reg, col_reg}<16'b0010100101100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100101100110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010100101100111) && ({row_reg, col_reg}<16'b0010100101101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010100101101001) && ({row_reg, col_reg}<16'b0010100101101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010100101101011) && ({row_reg, col_reg}<16'b0010100101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100101101110) && ({row_reg, col_reg}<16'b0010100101110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010100101110000) && ({row_reg, col_reg}<16'b0010100101110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100101110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100101110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100101110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100101110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100101110110) && ({row_reg, col_reg}<16'b0010100101111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010100101111000) && ({row_reg, col_reg}<16'b0010100101111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100101111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010100101111011) && ({row_reg, col_reg}<16'b0010100101111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100101111101) && ({row_reg, col_reg}<16'b0010100110000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010100110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100110000010) && ({row_reg, col_reg}<16'b0010100110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010100110010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100110010101) && ({row_reg, col_reg}<16'b0010100110011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100110011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010100110011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010100110011100) && ({row_reg, col_reg}<16'b0010100110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100110011111) && ({row_reg, col_reg}<16'b0010100110100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010100110100001) && ({row_reg, col_reg}<16'b0010100110100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100110100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100110100101) && ({row_reg, col_reg}<16'b0010100110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100110101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100110101001) && ({row_reg, col_reg}<16'b0010100110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100110101011) && ({row_reg, col_reg}<16'b0010100110101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010100110101110) && ({row_reg, col_reg}<16'b0010100110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010100110110000) && ({row_reg, col_reg}<16'b0010100110110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010100110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100110110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100110110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010100110110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010100110110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010100110111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010100110111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010100110111010) && ({row_reg, col_reg}<16'b0010100110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010100110111110) && ({row_reg, col_reg}<16'b0010100111000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100111000001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010100111000010) && ({row_reg, col_reg}<16'b0010100111000100)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}>=16'b0010100111000100) && ({row_reg, col_reg}<16'b0010100111001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010100111001000) && ({row_reg, col_reg}<16'b0010100111001010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010100111001010) && ({row_reg, col_reg}<16'b0010100111001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100111001110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010100111001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100111010000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0010100111010001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010100111010010)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0010100111010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100111010100) && ({row_reg, col_reg}<16'b0010100111010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100111010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010100111010111) && ({row_reg, col_reg}<16'b0010100111011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100111011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010100111011010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010100111011011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010100111011100) && ({row_reg, col_reg}<16'b0010100111011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100111011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010100111011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010100111100000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010100111100001)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0010100111100010) && ({row_reg, col_reg}<16'b0010100111100100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010100111100100) && ({row_reg, col_reg}<16'b0010100111100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100111100110) && ({row_reg, col_reg}<16'b0010100111101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010100111101010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010100111101011) && ({row_reg, col_reg}<16'b0010100111101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100111101101) && ({row_reg, col_reg}<16'b0010100111101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010100111101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010100111110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100111110001) && ({row_reg, col_reg}<16'b0010100111110011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010100111110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100111110100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010100111110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100111110110) && ({row_reg, col_reg}<16'b0010100111111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010100111111000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010100111111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010100111111010) && ({row_reg, col_reg}<16'b0010100111111100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010100111111100) && ({row_reg, col_reg}<16'b0010100111111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010100111111110)) color_data = 12'b001100110010;

		if(({row_reg, col_reg}==16'b0010100111111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010101000000000) && ({row_reg, col_reg}<16'b0010101000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101000000101) && ({row_reg, col_reg}<16'b0010101000000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101000000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010101000001000) && ({row_reg, col_reg}<16'b0010101000001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101000001011) && ({row_reg, col_reg}<16'b0010101000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101000010010) && ({row_reg, col_reg}<16'b0010101000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010101000011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101000011010) && ({row_reg, col_reg}<16'b0010101000100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101000100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101000100011) && ({row_reg, col_reg}<16'b0010101000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010101000101010) && ({row_reg, col_reg}<16'b0010101000110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101000110000) && ({row_reg, col_reg}<16'b0010101000110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101000110011) && ({row_reg, col_reg}<16'b0010101000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101000110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101000110110) && ({row_reg, col_reg}<16'b0010101000111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010101000111110) && ({row_reg, col_reg}<16'b0010101001000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101001000001) && ({row_reg, col_reg}<16'b0010101001000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101001000011) && ({row_reg, col_reg}<16'b0010101001000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101001000101) && ({row_reg, col_reg}<16'b0010101001001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101001001010) && ({row_reg, col_reg}<16'b0010101001001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101001001100) && ({row_reg, col_reg}<16'b0010101001010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010101001010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101001010100) && ({row_reg, col_reg}<16'b0010101001011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101001011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101001011110) && ({row_reg, col_reg}<16'b0010101001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010101001100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101001100010) && ({row_reg, col_reg}<16'b0010101001100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101001100100) && ({row_reg, col_reg}<16'b0010101001100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010101001100110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010101001100111) && ({row_reg, col_reg}<16'b0010101001101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101001101001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0010101001101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010101001101011) && ({row_reg, col_reg}<16'b0010101001101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101001101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101001101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010101001110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101001110001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0010101001110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010101001110011) && ({row_reg, col_reg}<16'b0010101001110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101001110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010101001111000) && ({row_reg, col_reg}<16'b0010101001111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101001111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010101001111011) && ({row_reg, col_reg}<16'b0010101001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101001111101) && ({row_reg, col_reg}<16'b0010101010000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101010000010) && ({row_reg, col_reg}<16'b0010101010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010101010010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101010010101) && ({row_reg, col_reg}<16'b0010101010011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101010011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010101010011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010101010011100) && ({row_reg, col_reg}<16'b0010101010100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101010100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101010100001) && ({row_reg, col_reg}<16'b0010101010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101010100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010101010100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101010100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010101010100110) && ({row_reg, col_reg}<16'b0010101010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101010101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101010101001) && ({row_reg, col_reg}<16'b0010101010101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101010101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010101010101100) && ({row_reg, col_reg}<16'b0010101010101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101010101110) && ({row_reg, col_reg}<16'b0010101010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101010110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010101010110001) && ({row_reg, col_reg}<16'b0010101010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101010110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010101010110110) && ({row_reg, col_reg}<16'b0010101010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101010111000) && ({row_reg, col_reg}<16'b0010101010111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101010111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010101010111100) && ({row_reg, col_reg}<16'b0010101010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010101010111110) && ({row_reg, col_reg}<16'b0010101011000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010101011000001) && ({row_reg, col_reg}<16'b0010101011000100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010101011000100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010101011000101) && ({row_reg, col_reg}<16'b0010101011001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010101011001000) && ({row_reg, col_reg}<16'b0010101011001010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010101011001010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010101011001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010101011001100) && ({row_reg, col_reg}<16'b0010101011001111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010101011001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101011010000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0010101011010001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010101011010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101011010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010101011010100) && ({row_reg, col_reg}<16'b0010101011010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101011010110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010101011010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010101011011000) && ({row_reg, col_reg}<16'b0010101011011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101011011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010101011011011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010101011011100) && ({row_reg, col_reg}<16'b0010101011011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101011011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010101011011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101011100000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010101011100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101011100010)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0010101011100011) && ({row_reg, col_reg}<16'b0010101011100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010101011100110) && ({row_reg, col_reg}<16'b0010101011101000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101011101000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0010101011101001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010101011101010) && ({row_reg, col_reg}<16'b0010101011101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101011101100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010101011101101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101011101110)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0010101011101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010101011110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101011110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101011110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010101011110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101011110100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101011110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010101011110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101011110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101011111000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0010101011111001) && ({row_reg, col_reg}<16'b0010101011111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101011111100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010101011111101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010101011111110)) color_data = 12'b001100110001;

		if(({row_reg, col_reg}==16'b0010101011111111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010101100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101100000001) && ({row_reg, col_reg}<16'b0010101100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101100000101) && ({row_reg, col_reg}<16'b0010101100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0010101100001000) && ({row_reg, col_reg}<16'b0010101100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101100001011) && ({row_reg, col_reg}<16'b0010101100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101100001111) && ({row_reg, col_reg}<16'b0010101100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101100010010) && ({row_reg, col_reg}<16'b0010101100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010101100011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101100011010) && ({row_reg, col_reg}<16'b0010101100100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101100100001) && ({row_reg, col_reg}<16'b0010101100100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101100100011) && ({row_reg, col_reg}<16'b0010101100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010101100101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101100101011) && ({row_reg, col_reg}<16'b0010101100110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101100110000) && ({row_reg, col_reg}<16'b0010101100110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101100110010) && ({row_reg, col_reg}<16'b0010101100110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101100110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101100110111) && ({row_reg, col_reg}<16'b0010101100111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010101100111110) && ({row_reg, col_reg}<16'b0010101101000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101101000001) && ({row_reg, col_reg}<16'b0010101101000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101101000100) && ({row_reg, col_reg}<16'b0010101101000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101101000110) && ({row_reg, col_reg}<16'b0010101101001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101101001010) && ({row_reg, col_reg}<16'b0010101101001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101101001100) && ({row_reg, col_reg}<16'b0010101101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010101101010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101101010100) && ({row_reg, col_reg}<16'b0010101101011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101101011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101101011110) && ({row_reg, col_reg}<16'b0010101101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010101101100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101101100010) && ({row_reg, col_reg}<16'b0010101101100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101101100100) && ({row_reg, col_reg}<16'b0010101101100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010101101100110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010101101100111) && ({row_reg, col_reg}<16'b0010101101101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101101101001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0010101101101010) && ({row_reg, col_reg}<16'b0010101101101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010101101101100) && ({row_reg, col_reg}<16'b0010101101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010101101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101101101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010101101110000) && ({row_reg, col_reg}<16'b0010101101110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101101110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010101101110011) && ({row_reg, col_reg}<16'b0010101101110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101101110111) && ({row_reg, col_reg}<16'b0010101101111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010101101111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010101101111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101101111011) && ({row_reg, col_reg}<16'b0010101101111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101101111101) && ({row_reg, col_reg}<16'b0010101110000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010101110000010) && ({row_reg, col_reg}<16'b0010101110010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010101110010101) && ({row_reg, col_reg}<16'b0010101110011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101110011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010101110011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010101110011100) && ({row_reg, col_reg}<16'b0010101110100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010101110100010) && ({row_reg, col_reg}<16'b0010101110100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010101110100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010101110100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101110100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010101110101000) && ({row_reg, col_reg}<16'b0010101110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101110110000) && ({row_reg, col_reg}<16'b0010101110110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010101110110010) && ({row_reg, col_reg}<16'b0010101110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010101110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010101110110110) && ({row_reg, col_reg}<16'b0010101110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010101110111000) && ({row_reg, col_reg}<16'b0010101110111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010101110111011) && ({row_reg, col_reg}<16'b0010101110111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010101110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010101110111110) && ({row_reg, col_reg}<16'b0010101111000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101111000001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010101111000010)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0010101111000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010101111000100) && ({row_reg, col_reg}<16'b0010101111000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010101111000111) && ({row_reg, col_reg}<16'b0010101111001011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010101111001011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010101111001100) && ({row_reg, col_reg}<16'b0010101111001111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010101111001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101111010000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0010101111010001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010101111010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101111010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010101111010100) && ({row_reg, col_reg}<16'b0010101111010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101111010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010101111010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010101111011000) && ({row_reg, col_reg}<16'b0010101111011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010101111011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010101111011011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010101111011100) && ({row_reg, col_reg}<16'b0010101111011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101111011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010101111011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010101111100000) && ({row_reg, col_reg}<16'b0010101111100010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101111100010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010101111100011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010101111100100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010101111100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010101111100110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010101111100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101111101000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0010101111101001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101111101010)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0010101111101011)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0010101111101100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010101111101101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0010101111101110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101111101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010101111110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101111110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101111110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010101111110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101111110100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010101111110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010101111110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010101111110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010101111111000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0010101111111001) && ({row_reg, col_reg}<16'b0010101111111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010101111111100) && ({row_reg, col_reg}<16'b0010101111111111)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}==16'b0010101111111111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010110000000000) && ({row_reg, col_reg}<16'b0010110000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110000000110) && ({row_reg, col_reg}<16'b0010110000001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110000001011) && ({row_reg, col_reg}<16'b0010110000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110000001111) && ({row_reg, col_reg}<16'b0010110000010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110000010010) && ({row_reg, col_reg}<16'b0010110000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110000011001) && ({row_reg, col_reg}<16'b0010110000011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110000011011) && ({row_reg, col_reg}<16'b0010110000100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110000100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110000100011) && ({row_reg, col_reg}<16'b0010110000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010110000101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110000101011) && ({row_reg, col_reg}<16'b0010110000110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110000110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110000110110) && ({row_reg, col_reg}<16'b0010110001000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010110001000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110001000001) && ({row_reg, col_reg}<16'b0010110001001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110001001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110001001100) && ({row_reg, col_reg}<16'b0010110001010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010110001010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110001010100) && ({row_reg, col_reg}<16'b0010110001011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110001011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110001011110) && ({row_reg, col_reg}<16'b0010110001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010110001100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010110001100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110001100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110001100100) && ({row_reg, col_reg}<16'b0010110001100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010110001100110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110001100111) && ({row_reg, col_reg}<16'b0010110001101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110001101001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0010110001101010) && ({row_reg, col_reg}<16'b0010110001101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010110001101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110001101101) && ({row_reg, col_reg}<16'b0010110001101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110001101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110001110000) && ({row_reg, col_reg}<16'b0010110001110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110001110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010110001110100) && ({row_reg, col_reg}<16'b0010110001110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110001110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110001110111) && ({row_reg, col_reg}<16'b0010110001111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010110001111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010110001111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110001111011) && ({row_reg, col_reg}<16'b0010110001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110001111101) && ({row_reg, col_reg}<16'b0010110010000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110010000010) && ({row_reg, col_reg}<16'b0010110010010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010110010010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110010010110) && ({row_reg, col_reg}<16'b0010110010011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110010011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010110010011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110010011100) && ({row_reg, col_reg}<16'b0010110010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110010100011) && ({row_reg, col_reg}<16'b0010110010100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110010100101) && ({row_reg, col_reg}<16'b0010110010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110010101000) && ({row_reg, col_reg}<16'b0010110010101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110010101011) && ({row_reg, col_reg}<16'b0010110010101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110010101101) && ({row_reg, col_reg}<16'b0010110010110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110010110001) && ({row_reg, col_reg}<16'b0010110010110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110010110011) && ({row_reg, col_reg}<16'b0010110010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110010110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010110010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110010110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110010111000) && ({row_reg, col_reg}<16'b0010110010111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010110010111011) && ({row_reg, col_reg}<16'b0010110010111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010110010111101) && ({row_reg, col_reg}<16'b0010110011000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110011000001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010110011000010)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0010110011000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010110011000100) && ({row_reg, col_reg}<16'b0010110011001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010110011001000) && ({row_reg, col_reg}<16'b0010110011001011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010110011001011) && ({row_reg, col_reg}<16'b0010110011001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110011001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010110011001110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010110011001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010110011010000) && ({row_reg, col_reg}<16'b0010110011010011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010110011010011) && ({row_reg, col_reg}<16'b0010110011010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110011010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110011011000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010110011011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110011011010) && ({row_reg, col_reg}<16'b0010110011011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010110011011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010110011011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010110011011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110011011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010110011100000) && ({row_reg, col_reg}<16'b0010110011100010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010110011100010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010110011100011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010110011100100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010110011100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010110011100110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010110011100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010110011101000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0010110011101001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010110011101010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010110011101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010110011101100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0010110011101101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010110011101110)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0010110011101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110011110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010110011110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110011110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010110011110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110011110100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010110011110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110011110110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010110011110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110011111000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0010110011111001) && ({row_reg, col_reg}<16'b0010110011111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110011111100)) color_data = 12'b001100110010;

		if(({row_reg, col_reg}>=16'b0010110011111101) && ({row_reg, col_reg}<16'b0010110100000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010110100000000) && ({row_reg, col_reg}<16'b0010110100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110100000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010110100000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110100000111) && ({row_reg, col_reg}<16'b0010110100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110100001101) && ({row_reg, col_reg}<16'b0010110100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110100001111) && ({row_reg, col_reg}<16'b0010110100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110100010010) && ({row_reg, col_reg}<16'b0010110100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110100011010) && ({row_reg, col_reg}<16'b0010110100011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010110100011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110100011101) && ({row_reg, col_reg}<16'b0010110100011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110100011111) && ({row_reg, col_reg}<16'b0010110100100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110100100001) && ({row_reg, col_reg}<16'b0010110100100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110100100011) && ({row_reg, col_reg}<16'b0010110100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010110100101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110100101011) && ({row_reg, col_reg}<16'b0010110100110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110100110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110100110101) && ({row_reg, col_reg}<16'b0010110100111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110100111011) && ({row_reg, col_reg}<16'b0010110100111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110100111101) && ({row_reg, col_reg}<16'b0010110101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110101000001) && ({row_reg, col_reg}<16'b0010110101000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110101000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110101000100) && ({row_reg, col_reg}<16'b0010110101000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110101000110) && ({row_reg, col_reg}<16'b0010110101001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010110101001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110101001010) && ({row_reg, col_reg}<16'b0010110101001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110101001100) && ({row_reg, col_reg}<16'b0010110101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010110101010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110101010100) && ({row_reg, col_reg}<16'b0010110101010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110101010110) && ({row_reg, col_reg}<16'b0010110101011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010110101011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110101011011) && ({row_reg, col_reg}<16'b0010110101011110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110101011110) && ({row_reg, col_reg}<16'b0010110101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010110101100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110101100010) && ({row_reg, col_reg}<16'b0010110101100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110101100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010110101100110) && ({row_reg, col_reg}<16'b0010110101101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110101101000) && ({row_reg, col_reg}<16'b0010110101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010110101101010) && ({row_reg, col_reg}<16'b0010110101101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010110101101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110101101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110101110000) && ({row_reg, col_reg}<16'b0010110101110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010110101110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110101110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010110101110100) && ({row_reg, col_reg}<16'b0010110101110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110101110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010110101111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010110101111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110101111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110101111011) && ({row_reg, col_reg}<16'b0010110101111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110101111101) && ({row_reg, col_reg}<16'b0010110101111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110101111111) && ({row_reg, col_reg}<16'b0010110110000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110110000010) && ({row_reg, col_reg}<16'b0010110110010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110110010110) && ({row_reg, col_reg}<16'b0010110110011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010110110011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010110110011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110110011100) && ({row_reg, col_reg}<16'b0010110110100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110110100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010110110100001) && ({row_reg, col_reg}<16'b0010110110100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110110100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110110100100) && ({row_reg, col_reg}<16'b0010110110100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110110100110) && ({row_reg, col_reg}<16'b0010110110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010110110101000) && ({row_reg, col_reg}<16'b0010110110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010110110101011) && ({row_reg, col_reg}<16'b0010110110101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010110110101101) && ({row_reg, col_reg}<16'b0010110110110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010110110110011) && ({row_reg, col_reg}<16'b0010110110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110110110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010110110110110) && ({row_reg, col_reg}<16'b0010110110111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010110110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010110110111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010110110111011) && ({row_reg, col_reg}<16'b0010110110111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010110110111101) && ({row_reg, col_reg}<16'b0010110110111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110110111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010110111000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110111000001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010110111000010)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0010110111000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010110111000100) && ({row_reg, col_reg}<16'b0010110111001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010110111001001) && ({row_reg, col_reg}<16'b0010110111001100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010110111001100) && ({row_reg, col_reg}<16'b0010110111001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110111001110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010110111001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110111010000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010110111010001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010110111010010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010110111010011) && ({row_reg, col_reg}<16'b0010110111010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110111010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110111011000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010110111011001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010110111011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010110111011011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010110111011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010110111011101) && ({row_reg, col_reg}<16'b0010110111011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110111011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010110111100000) && ({row_reg, col_reg}<16'b0010110111100010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010110111100010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010110111100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010110111100100) && ({row_reg, col_reg}<16'b0010110111100110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0010110111100110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010110111100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010110111101000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0010110111101001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0010110111101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010110111101011) && ({row_reg, col_reg}<16'b0010110111101110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010110111101110)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0010110111101111) && ({row_reg, col_reg}<16'b0010110111110001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010110111110001)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010110111110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010110111110011) && ({row_reg, col_reg}<16'b0010110111110101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010110111110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010110111110110) && ({row_reg, col_reg}<16'b0010110111111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010110111111000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0010110111111001) && ({row_reg, col_reg}<16'b0010110111111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010110111111100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010110111111101)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010110111111110)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}==16'b0010110111111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111000000000) && ({row_reg, col_reg}<16'b0010111000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111000000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111000000110) && ({row_reg, col_reg}<16'b0010111000001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010111000001000) && ({row_reg, col_reg}<16'b0010111000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111000001100) && ({row_reg, col_reg}<16'b0010111000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111000001111) && ({row_reg, col_reg}<16'b0010111000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111000010010) && ({row_reg, col_reg}<16'b0010111000011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010111000011010) && ({row_reg, col_reg}<16'b0010111000100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111000100010) && ({row_reg, col_reg}<16'b0010111000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010111000101010) && ({row_reg, col_reg}<16'b0010111000110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111000110101) && ({row_reg, col_reg}<16'b0010111000111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010111000111010) && ({row_reg, col_reg}<16'b0010111000111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111000111101) && ({row_reg, col_reg}<16'b0010111001000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010111001000001) && ({row_reg, col_reg}<16'b0010111001001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111001001011) && ({row_reg, col_reg}<16'b0010111001010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010111001010100) && ({row_reg, col_reg}<16'b0010111001011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111001011100) && ({row_reg, col_reg}<16'b0010111001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010111001100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111001100010) && ({row_reg, col_reg}<16'b0010111001100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111001100101) && ({row_reg, col_reg}<16'b0010111001100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010111001100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010111001101000) && ({row_reg, col_reg}<16'b0010111001101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111001101010) && ({row_reg, col_reg}<16'b0010111001101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111001101100) && ({row_reg, col_reg}<16'b0010111001101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111001101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111001101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111001110000) && ({row_reg, col_reg}<16'b0010111001110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010111001110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010111001110011) && ({row_reg, col_reg}<16'b0010111001110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111001110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111001111000) && ({row_reg, col_reg}<16'b0010111001111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111001111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010111001111011) && ({row_reg, col_reg}<16'b0010111001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111001111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111001111110) && ({row_reg, col_reg}<16'b0010111010000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010111010000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111010000010) && ({row_reg, col_reg}<16'b0010111010010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010111010010011) && ({row_reg, col_reg}<16'b0010111010010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010111010010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010111010010110) && ({row_reg, col_reg}<16'b0010111010011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111010011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010111010011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010111010011100) && ({row_reg, col_reg}<16'b0010111010100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111010100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111010100001) && ({row_reg, col_reg}<16'b0010111010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111010100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111010100100) && ({row_reg, col_reg}<16'b0010111010100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111010100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111010100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010111010101000) && ({row_reg, col_reg}<16'b0010111010101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111010101011) && ({row_reg, col_reg}<16'b0010111010101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010111010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111010101110) && ({row_reg, col_reg}<16'b0010111010110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111010110011) && ({row_reg, col_reg}<16'b0010111010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111010110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010111010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111010110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010111010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111010111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111010111011) && ({row_reg, col_reg}<16'b0010111010111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111010111101) && ({row_reg, col_reg}<16'b0010111010111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111010111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010111011000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111011000001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0010111011000010)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0010111011000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010111011000100) && ({row_reg, col_reg}<16'b0010111011001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111011001010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010111011001011) && ({row_reg, col_reg}<16'b0010111011001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111011001101)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0010111011001110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010111011001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010111011010000) && ({row_reg, col_reg}<16'b0010111011010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010111011010010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0010111011010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111011010100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010111011010101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0010111011010110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0010111011010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010111011011000) && ({row_reg, col_reg}<16'b0010111011011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111011011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010111011011011) && ({row_reg, col_reg}<16'b0010111011011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010111011011101) && ({row_reg, col_reg}<16'b0010111011100000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010111011100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111011100001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010111011100010) && ({row_reg, col_reg}<16'b0010111011100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111011100110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010111011100111) && ({row_reg, col_reg}<16'b0010111011101011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010111011101011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111011101100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010111011101101)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}>=16'b0010111011101110) && ({row_reg, col_reg}<16'b0010111011110000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0010111011110000) && ({row_reg, col_reg}<16'b0010111011110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010111011110010)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0010111011110011) && ({row_reg, col_reg}<16'b0010111011110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010111011110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010111011110110) && ({row_reg, col_reg}<16'b0010111011111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111011111000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010111011111001) && ({row_reg, col_reg}<16'b0010111011111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010111011111101) && ({row_reg, col_reg}<16'b0010111011111111)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}==16'b0010111011111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111100000000) && ({row_reg, col_reg}<16'b0010111100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111100000110) && ({row_reg, col_reg}<16'b0010111100001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010111100001000) && ({row_reg, col_reg}<16'b0010111100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0010111100001101) && ({row_reg, col_reg}<16'b0010111100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111100010001) && ({row_reg, col_reg}<16'b0010111100111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010111100111010) && ({row_reg, col_reg}<16'b0010111100111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111100111101) && ({row_reg, col_reg}<16'b0010111101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010111101100001) && ({row_reg, col_reg}<16'b0010111101100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111101100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010111101100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111101100110) && ({row_reg, col_reg}<16'b0010111101101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111101101000) && ({row_reg, col_reg}<16'b0010111101101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111101101010) && ({row_reg, col_reg}<16'b0010111101101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111101101100) && ({row_reg, col_reg}<16'b0010111101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111101101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111101110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010111101110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111101110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010111101110011) && ({row_reg, col_reg}<16'b0010111101110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111101110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111101111000) && ({row_reg, col_reg}<16'b0010111101111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111101111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010111101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111101111100) && ({row_reg, col_reg}<16'b0010111101111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010111101111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111101111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010111110000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0010111110000010) && ({row_reg, col_reg}<16'b0010111110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0010111110010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010111110010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111110010110) && ({row_reg, col_reg}<16'b0010111110011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111110011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111110011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010111110011100) && ({row_reg, col_reg}<16'b0010111110100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111110100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0010111110100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111110100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111110100011) && ({row_reg, col_reg}<16'b0010111110100110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010111110100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0010111110100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0010111110101000) && ({row_reg, col_reg}<16'b0010111110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111110101011) && ({row_reg, col_reg}<16'b0010111110101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010111110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0010111110101110) && ({row_reg, col_reg}<16'b0010111110110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0010111110110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0010111110110100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0010111110110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010111110110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0010111110110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0010111110111000) && ({row_reg, col_reg}<16'b0010111110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111110111010) && ({row_reg, col_reg}<16'b0010111110111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0010111110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111110111110) && ({row_reg, col_reg}<16'b0010111111000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111111000000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0010111111000001) && ({row_reg, col_reg}<16'b0010111111000100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010111111000100) && ({row_reg, col_reg}<16'b0010111111000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0010111111000110) && ({row_reg, col_reg}<16'b0010111111001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010111111001001) && ({row_reg, col_reg}<16'b0010111111001011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010111111001011) && ({row_reg, col_reg}<16'b0010111111001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111111001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111111001111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0010111111010000) && ({row_reg, col_reg}<16'b0010111111010011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010111111010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111111010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010111111010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111111010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0010111111010111) && ({row_reg, col_reg}<16'b0010111111011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0010111111011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0010111111011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0010111111011011) && ({row_reg, col_reg}<16'b0010111111011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0010111111011110) && ({row_reg, col_reg}<16'b0010111111100000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010111111100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111111100001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010111111100010) && ({row_reg, col_reg}<16'b0010111111100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111111100101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0010111111100110) && ({row_reg, col_reg}<16'b0010111111101000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010111111101000) && ({row_reg, col_reg}<16'b0010111111101010)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0010111111101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0010111111101011) && ({row_reg, col_reg}<16'b0010111111101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111111101101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0010111111101110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0010111111101111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0010111111110000) && ({row_reg, col_reg}<16'b0010111111110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0010111111110010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0010111111110011) && ({row_reg, col_reg}<16'b0010111111110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0010111111110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0010111111110110) && ({row_reg, col_reg}<16'b0010111111111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0010111111111000) && ({row_reg, col_reg}<16'b0010111111111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0010111111111110)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}==16'b0010111111111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011000000000000) && ({row_reg, col_reg}<16'b0011000000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000000000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000000000110) && ({row_reg, col_reg}<16'b0011000000001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011000000001000) && ({row_reg, col_reg}<16'b0011000000001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000000001011) && ({row_reg, col_reg}<16'b0011000000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000000010010) && ({row_reg, col_reg}<16'b0011000000111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011000000111010) && ({row_reg, col_reg}<16'b0011000000111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011000000111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000000111101) && ({row_reg, col_reg}<16'b0011000001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011000001100001) && ({row_reg, col_reg}<16'b0011000001100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000001100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011000001100100) && ({row_reg, col_reg}<16'b0011000001100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000001100111) && ({row_reg, col_reg}<16'b0011000001101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011000001101101) && ({row_reg, col_reg}<16'b0011000001101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000001101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011000001110000) && ({row_reg, col_reg}<16'b0011000001110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000001110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011000001110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000001110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011000001110101) && ({row_reg, col_reg}<16'b0011000001110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000001110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011000001111000) && ({row_reg, col_reg}<16'b0011000001111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000001111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011000001111011) && ({row_reg, col_reg}<16'b0011000001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000001111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011000001111110) && ({row_reg, col_reg}<16'b0011000010000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011000010000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011000010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000010000010) && ({row_reg, col_reg}<16'b0011000010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011000010010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000010010101) && ({row_reg, col_reg}<16'b0011000010010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000010010111) && ({row_reg, col_reg}<16'b0011000010011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011000010011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011000010011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011000010011100) && ({row_reg, col_reg}<16'b0011000010100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000010100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011000010100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000010100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000010100011) && ({row_reg, col_reg}<16'b0011000010100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011000010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000010100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011000010100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011000010101000) && ({row_reg, col_reg}<16'b0011000010101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000010101011) && ({row_reg, col_reg}<16'b0011000010101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011000010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000010101110) && ({row_reg, col_reg}<16'b0011000010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000010110000) && ({row_reg, col_reg}<16'b0011000010110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011000010110011) && ({row_reg, col_reg}<16'b0011000010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000010110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011000010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000010110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011000010111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011000010111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011000010111011) && ({row_reg, col_reg}<16'b0011000010111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011000010111101) && ({row_reg, col_reg}<16'b0011000010111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000010111111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011000011000000) && ({row_reg, col_reg}<16'b0011000011000100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011000011000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011000011000101) && ({row_reg, col_reg}<16'b0011000011001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011000011001001) && ({row_reg, col_reg}<16'b0011000011001011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011000011001011) && ({row_reg, col_reg}<16'b0011000011001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000011001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000011001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011000011010000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0011000011010001) && ({row_reg, col_reg}<16'b0011000011010011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011000011010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011000011010100) && ({row_reg, col_reg}<16'b0011000011010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011000011010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011000011010111) && ({row_reg, col_reg}<16'b0011000011011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011000011011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011000011011010) && ({row_reg, col_reg}<16'b0011000011011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011000011011100) && ({row_reg, col_reg}<16'b0011000011011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000011011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011000011100000)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0011000011100001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0011000011100010) && ({row_reg, col_reg}<16'b0011000011100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000011100100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0011000011100101) && ({row_reg, col_reg}<16'b0011000011100111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011000011100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011000011101000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0011000011101001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011000011101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011000011101011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000011101100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011000011101101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0011000011101110) && ({row_reg, col_reg}<16'b0011000011110000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011000011110000) && ({row_reg, col_reg}<16'b0011000011110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011000011110010)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0011000011110011) && ({row_reg, col_reg}<16'b0011000011110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011000011110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011000011110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000011110111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011000011111000) && ({row_reg, col_reg}<16'b0011000011111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000011111010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011000011111011) && ({row_reg, col_reg}<16'b0011000011111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000011111110)) color_data = 12'b010000100001;

		if(({row_reg, col_reg}==16'b0011000011111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011000100000000) && ({row_reg, col_reg}<16'b0011000100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000100000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000100000111) && ({row_reg, col_reg}<16'b0011000100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011000100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000100001010) && ({row_reg, col_reg}<16'b0011000100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000100010001) && ({row_reg, col_reg}<16'b0011000100111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011000100111011) && ({row_reg, col_reg}<16'b0011000100111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000100111110) && ({row_reg, col_reg}<16'b0011000101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011000101100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000101100010) && ({row_reg, col_reg}<16'b0011000101101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000101101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011000101101101) && ({row_reg, col_reg}<16'b0011000101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000101110000) && ({row_reg, col_reg}<16'b0011000101110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011000101110011) && ({row_reg, col_reg}<16'b0011000101110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000101110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011000101111000) && ({row_reg, col_reg}<16'b0011000101111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011000101111011) && ({row_reg, col_reg}<16'b0011000101111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000101111101) && ({row_reg, col_reg}<16'b0011000110000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011000110000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011000110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000110000010) && ({row_reg, col_reg}<16'b0011000110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011000110010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011000110010101) && ({row_reg, col_reg}<16'b0011000110011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000110011000) && ({row_reg, col_reg}<16'b0011000110011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000110011010) && ({row_reg, col_reg}<16'b0011000110011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011000110011100) && ({row_reg, col_reg}<16'b0011000110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000110011111) && ({row_reg, col_reg}<16'b0011000110100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011000110100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000110100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000110100011) && ({row_reg, col_reg}<16'b0011000110100110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011000110100110) && ({row_reg, col_reg}<16'b0011000110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000110101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011000110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000110101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011000110101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011000110101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011000110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011000110101110) && ({row_reg, col_reg}<16'b0011000110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011000110110000) && ({row_reg, col_reg}<16'b0011000110110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011000110110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011000110110011) && ({row_reg, col_reg}<16'b0011000110110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011000110110110) && ({row_reg, col_reg}<16'b0011000110111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011000110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011000110111001) && ({row_reg, col_reg}<16'b0011000110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000110111011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0011000110111100) && ({row_reg, col_reg}<16'b0011000110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011000110111110) && ({row_reg, col_reg}<16'b0011000111000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011000111000010) && ({row_reg, col_reg}<16'b0011000111000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011000111000101) && ({row_reg, col_reg}<16'b0011000111001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011000111001000) && ({row_reg, col_reg}<16'b0011000111001010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011000111001010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011000111001011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011000111001100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011000111001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011000111001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000111001111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0011000111010000) && ({row_reg, col_reg}<16'b0011000111010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011000111010010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0011000111010011) && ({row_reg, col_reg}<16'b0011000111010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000111010110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011000111010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011000111011000) && ({row_reg, col_reg}<16'b0011000111011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011000111011100) && ({row_reg, col_reg}<16'b0011000111100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000111100000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0011000111100001) && ({row_reg, col_reg}<16'b0011000111100011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0011000111100011) && ({row_reg, col_reg}<16'b0011000111100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000111100101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011000111100110) && ({row_reg, col_reg}<16'b0011000111101000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011000111101000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0011000111101001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0011000111101010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0011000111101011) && ({row_reg, col_reg}<16'b0011000111101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000111101101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011000111101110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011000111101111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011000111110000) && ({row_reg, col_reg}<16'b0011000111110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011000111110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011000111110011) && ({row_reg, col_reg}<16'b0011000111110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011000111110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000111110110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011000111110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011000111111000) && ({row_reg, col_reg}<16'b0011000111111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000111111010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011000111111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000111111100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011000111111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011000111111110)) color_data = 12'b010000100001;

		if(({row_reg, col_reg}==16'b0011000111111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011001000000000) && ({row_reg, col_reg}<16'b0011001000000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001000000100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011001000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001000000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001000000111) && ({row_reg, col_reg}<16'b0011001000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011001000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011001000001010) && ({row_reg, col_reg}<16'b0011001000001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011001000001100) && ({row_reg, col_reg}<16'b0011001000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001000010010) && ({row_reg, col_reg}<16'b0011001000111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011001000111100) && ({row_reg, col_reg}<16'b0011001000111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001000111110) && ({row_reg, col_reg}<16'b0011001001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011001001100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001001100010) && ({row_reg, col_reg}<16'b0011001001100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001001100100) && ({row_reg, col_reg}<16'b0011001001100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001001100110) && ({row_reg, col_reg}<16'b0011001001101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001001101000) && ({row_reg, col_reg}<16'b0011001001101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001001101010) && ({row_reg, col_reg}<16'b0011001001101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001001101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011001001101101) && ({row_reg, col_reg}<16'b0011001001110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001001110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011001001110110) && ({row_reg, col_reg}<16'b0011001001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001001111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011001001111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011001001111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011001001111011) && ({row_reg, col_reg}<16'b0011001001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001001111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001001111110) && ({row_reg, col_reg}<16'b0011001010000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011001010000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011001010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001010000010) && ({row_reg, col_reg}<16'b0011001010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011001010010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001010010101) && ({row_reg, col_reg}<16'b0011001010011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001010011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011001010011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001010011010) && ({row_reg, col_reg}<16'b0011001010011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011001010011100) && ({row_reg, col_reg}<16'b0011001010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001010011111) && ({row_reg, col_reg}<16'b0011001010100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001010100001) && ({row_reg, col_reg}<16'b0011001010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001010100011) && ({row_reg, col_reg}<16'b0011001010100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011001010100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011001010100110) && ({row_reg, col_reg}<16'b0011001010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011001010101000) && ({row_reg, col_reg}<16'b0011001010101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011001010101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011001010101100) && ({row_reg, col_reg}<16'b0011001010101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011001010101110) && ({row_reg, col_reg}<16'b0011001010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001010110000) && ({row_reg, col_reg}<16'b0011001010110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011001010110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011001010110011) && ({row_reg, col_reg}<16'b0011001010110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011001010110110) && ({row_reg, col_reg}<16'b0011001010111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011001010111000) && ({row_reg, col_reg}<16'b0011001010111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011001010111011) && ({row_reg, col_reg}<16'b0011001010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011001010111110) && ({row_reg, col_reg}<16'b0011001011000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001011000011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011001011000100) && ({row_reg, col_reg}<16'b0011001011000110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011001011000110) && ({row_reg, col_reg}<16'b0011001011001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001011001000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011001011001001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011001011001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001011001011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011001011001100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011001011001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001011001110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011001011001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011001011010000) && ({row_reg, col_reg}<16'b0011001011010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011001011010010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0011001011010011) && ({row_reg, col_reg}<16'b0011001011010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001011010101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011001011010110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011001011010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001011011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011001011011001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011001011011010) && ({row_reg, col_reg}<16'b0011001011011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011001011011100) && ({row_reg, col_reg}<16'b0011001011100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011001011100001) && ({row_reg, col_reg}<16'b0011001011100011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0011001011100011) && ({row_reg, col_reg}<16'b0011001011100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001011100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011001011100110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0011001011100111) && ({row_reg, col_reg}<16'b0011001011101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011001011101010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011001011101011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001011101100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011001011101101) && ({row_reg, col_reg}<16'b0011001011101111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011001011101111)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0011001011110000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011001011110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001011110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011001011110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001011110100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011001011110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001011110110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011001011110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001011111000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011001011111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001011111010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011001011111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001011111100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011001011111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001011111110)) color_data = 12'b010000100001;

		if(({row_reg, col_reg}==16'b0011001011111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011001100000000) && ({row_reg, col_reg}<16'b0011001100000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001100000100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011001100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001100000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011001100000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011001100001000) && ({row_reg, col_reg}<16'b0011001100001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011001100001010) && ({row_reg, col_reg}<16'b0011001100001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011001100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001100001101) && ({row_reg, col_reg}<16'b0011001100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001100010010) && ({row_reg, col_reg}<16'b0011001101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011001101100001) && ({row_reg, col_reg}<16'b0011001101100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001101100100) && ({row_reg, col_reg}<16'b0011001101100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001101100110) && ({row_reg, col_reg}<16'b0011001101101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001101101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001101101001) && ({row_reg, col_reg}<16'b0011001101101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001101101111) && ({row_reg, col_reg}<16'b0011001101110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001101110010) && ({row_reg, col_reg}<16'b0011001101110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001101110100) && ({row_reg, col_reg}<16'b0011001101110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011001101110110) && ({row_reg, col_reg}<16'b0011001101111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001101111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011001101111010) && ({row_reg, col_reg}<16'b0011001101111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001101111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011001101111111) && ({row_reg, col_reg}<16'b0011001110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001110000010) && ({row_reg, col_reg}<16'b0011001110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011001110010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001110010101) && ({row_reg, col_reg}<16'b0011001110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001110010111) && ({row_reg, col_reg}<16'b0011001110011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001110011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001110011010) && ({row_reg, col_reg}<16'b0011001110011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011001110011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011001110011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001110011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011001110011111) && ({row_reg, col_reg}<16'b0011001110100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011001110100001) && ({row_reg, col_reg}<16'b0011001110100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001110100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011001110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011001110100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011001110100110) && ({row_reg, col_reg}<16'b0011001110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011001110101000) && ({row_reg, col_reg}<16'b0011001110101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011001110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011001110101110) && ({row_reg, col_reg}<16'b0011001110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011001110110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011001110110001) && ({row_reg, col_reg}<16'b0011001110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011001110110011) && ({row_reg, col_reg}<16'b0011001110110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011001110110110) && ({row_reg, col_reg}<16'b0011001110111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011001110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011001110111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011001110111011) && ({row_reg, col_reg}<16'b0011001110111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011001110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011001110111110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001110111111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011001111000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001111000001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011001111000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011001111000011) && ({row_reg, col_reg}<16'b0011001111000110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011001111000110) && ({row_reg, col_reg}<16'b0011001111001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001111001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011001111001001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011001111001010) && ({row_reg, col_reg}<16'b0011001111001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011001111001110) && ({row_reg, col_reg}<16'b0011001111010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001111010000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011001111010001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011001111010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011001111010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001111010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011001111010101) && ({row_reg, col_reg}<16'b0011001111011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001111011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001111011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011001111011010) && ({row_reg, col_reg}<16'b0011001111011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011001111011100) && ({row_reg, col_reg}<16'b0011001111011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001111011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011001111100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011001111100001) && ({row_reg, col_reg}<16'b0011001111100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0011001111100101) && ({row_reg, col_reg}<16'b0011001111100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011001111100111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0011001111101000) && ({row_reg, col_reg}<16'b0011001111101011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0011001111101011) && ({row_reg, col_reg}<16'b0011001111101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001111101110)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0011001111101111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011001111110000) && ({row_reg, col_reg}<16'b0011001111110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001111110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001111110100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011001111110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001111110110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011001111110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001111111000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011001111111001) && ({row_reg, col_reg}<16'b0011001111111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011001111111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011001111111100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011001111111101)) color_data = 12'b010100110010;

		if(({row_reg, col_reg}>=16'b0011001111111110) && ({row_reg, col_reg}<16'b0011010000000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011010000000000) && ({row_reg, col_reg}<16'b0011010000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010000000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011010000000111) && ({row_reg, col_reg}<16'b0011010000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011010000001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010000001011) && ({row_reg, col_reg}<16'b0011010000001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011010000001101) && ({row_reg, col_reg}<16'b0011010000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010000010010) && ({row_reg, col_reg}<16'b0011010001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011010001100001) && ({row_reg, col_reg}<16'b0011010001100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010001100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011010001100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010001100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010001100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010001100111) && ({row_reg, col_reg}<16'b0011010001101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010001101001) && ({row_reg, col_reg}<16'b0011010001101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010001101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010001110000) && ({row_reg, col_reg}<16'b0011010001110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011010001110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010001110011) && ({row_reg, col_reg}<16'b0011010010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010010000010) && ({row_reg, col_reg}<16'b0011010010010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011010010010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011010010010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010010010101) && ({row_reg, col_reg}<16'b0011010010010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011010010010111) && ({row_reg, col_reg}<16'b0011010010011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010010011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010010011010) && ({row_reg, col_reg}<16'b0011010010011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011010010011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011010010011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010010011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010010100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010010100001) && ({row_reg, col_reg}<16'b0011010010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010010100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011010010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010010100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011010010100110) && ({row_reg, col_reg}<16'b0011010010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010010101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011010010101001) && ({row_reg, col_reg}<16'b0011010010101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010010101011) && ({row_reg, col_reg}<16'b0011010010101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011010010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010010101110) && ({row_reg, col_reg}<16'b0011010010110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010010110001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011010010110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011010010110011) && ({row_reg, col_reg}<16'b0011010010110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011010010110110) && ({row_reg, col_reg}<16'b0011010010111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011010010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011010010111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011010010111011) && ({row_reg, col_reg}<16'b0011010010111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011010010111101) && ({row_reg, col_reg}<16'b0011010010111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011010010111111) && ({row_reg, col_reg}<16'b0011010011000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011010011000001) && ({row_reg, col_reg}<16'b0011010011000011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0011010011000011) && ({row_reg, col_reg}<16'b0011010011000110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011010011000110) && ({row_reg, col_reg}<16'b0011010011001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011010011001000) && ({row_reg, col_reg}<16'b0011010011001010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011010011001010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0011010011001011) && ({row_reg, col_reg}<16'b0011010011001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010011001110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011010011001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010011010000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0011010011010001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011010011010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011010011010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011010011010100) && ({row_reg, col_reg}<16'b0011010011010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010011010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011010011010111) && ({row_reg, col_reg}<16'b0011010011011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010011011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011010011011010) && ({row_reg, col_reg}<16'b0011010011011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011010011011100) && ({row_reg, col_reg}<16'b0011010011011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010011011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010011011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011010011100000) && ({row_reg, col_reg}<16'b0011010011100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010011100100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0011010011100101) && ({row_reg, col_reg}<16'b0011010011100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011010011100111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011010011101000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0011010011101001) && ({row_reg, col_reg}<16'b0011010011101011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011010011101011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011010011101100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011010011101101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0011010011101110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011010011101111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0011010011110000) && ({row_reg, col_reg}<16'b0011010011110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010011110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010011110100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0011010011110101) && ({row_reg, col_reg}<16'b0011010011110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011010011110111) && ({row_reg, col_reg}<16'b0011010011111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010011111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010011111100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011010011111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010011111110)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}==16'b0011010011111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011010100000000) && ({row_reg, col_reg}<16'b0011010100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010100000101) && ({row_reg, col_reg}<16'b0011010100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011010100001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011010100001001) && ({row_reg, col_reg}<16'b0011010100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011010100001100) && ({row_reg, col_reg}<16'b0011010100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010100010010) && ({row_reg, col_reg}<16'b0011010101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011010101100001) && ({row_reg, col_reg}<16'b0011010101100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010101100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011010101100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010101100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010101100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010101100111) && ({row_reg, col_reg}<16'b0011010101101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010101101001) && ({row_reg, col_reg}<16'b0011010101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010101101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011010101101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010101110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011010101110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011010101110010) && ({row_reg, col_reg}<16'b0011010101110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011010101110101) && ({row_reg, col_reg}<16'b0011010101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010101111000) && ({row_reg, col_reg}<16'b0011010101111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010101111011) && ({row_reg, col_reg}<16'b0011010101111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011010101111101) && ({row_reg, col_reg}<16'b0011010110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010110000010) && ({row_reg, col_reg}<16'b0011010110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011010110010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010110010101) && ({row_reg, col_reg}<16'b0011010110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011010110010111) && ({row_reg, col_reg}<16'b0011010110011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010110011010) && ({row_reg, col_reg}<16'b0011010110011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010110011100) && ({row_reg, col_reg}<16'b0011010110100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010110100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011010110100001) && ({row_reg, col_reg}<16'b0011010110100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010110100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011010110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011010110100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010110100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011010110100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011010110101000) && ({row_reg, col_reg}<16'b0011010110101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010110101011) && ({row_reg, col_reg}<16'b0011010110101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011010110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011010110101110) && ({row_reg, col_reg}<16'b0011010110110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010110110001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011010110110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011010110110011) && ({row_reg, col_reg}<16'b0011010110110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011010110110110) && ({row_reg, col_reg}<16'b0011010110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011010110111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011010110111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011010110111011) && ({row_reg, col_reg}<16'b0011010110111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011010110111101) && ({row_reg, col_reg}<16'b0011010110111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011010110111111) && ({row_reg, col_reg}<16'b0011010111000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011010111000010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0011010111000011) && ({row_reg, col_reg}<16'b0011010111000110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011010111000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011010111000111) && ({row_reg, col_reg}<16'b0011010111001010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011010111001010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010111001011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011010111001100) && ({row_reg, col_reg}<16'b0011010111001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010111001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011010111001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010111010000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0011010111010001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011010111010010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011010111010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011010111010100) && ({row_reg, col_reg}<16'b0011010111010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011010111010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010111010111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011010111011000) && ({row_reg, col_reg}<16'b0011010111011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011010111011010) && ({row_reg, col_reg}<16'b0011010111011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011010111011100) && ({row_reg, col_reg}<16'b0011010111011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010111011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011010111011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010111100000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011010111100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0011010111100010) && ({row_reg, col_reg}<16'b0011010111100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011010111100100) && ({row_reg, col_reg}<16'b0011010111101000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0011010111101000) && ({row_reg, col_reg}<16'b0011010111101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011010111101010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011010111101011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0011010111101100) && ({row_reg, col_reg}<16'b0011010111101111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011010111101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010111110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011010111110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010111110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0011010111110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010111110100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011010111110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011010111110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011010111110111) && ({row_reg, col_reg}<16'b0011010111111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011010111111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011010111111100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011010111111101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011010111111110)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}==16'b0011010111111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011000000001) && ({row_reg, col_reg}<16'b0011011000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011000000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011000000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011011000000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011011000001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011011000001001) && ({row_reg, col_reg}<16'b0011011000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011000001100) && ({row_reg, col_reg}<16'b0011011000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011000010001) && ({row_reg, col_reg}<16'b0011011001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011011001100001) && ({row_reg, col_reg}<16'b0011011001100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011001100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011001100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011001100111) && ({row_reg, col_reg}<16'b0011011001101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011001101001) && ({row_reg, col_reg}<16'b0011011001101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011001101011) && ({row_reg, col_reg}<16'b0011011001101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011001101101) && ({row_reg, col_reg}<16'b0011011001110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011001110011) && ({row_reg, col_reg}<16'b0011011001110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011001110110) && ({row_reg, col_reg}<16'b0011011001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011001111000) && ({row_reg, col_reg}<16'b0011011001111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011001111011) && ({row_reg, col_reg}<16'b0011011001111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011001111110) && ({row_reg, col_reg}<16'b0011011010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011010000001) && ({row_reg, col_reg}<16'b0011011010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011011010010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011010010101) && ({row_reg, col_reg}<16'b0011011010010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011010010111) && ({row_reg, col_reg}<16'b0011011010011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011010011001) && ({row_reg, col_reg}<16'b0011011010011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011010011100) && ({row_reg, col_reg}<16'b0011011010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011010100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011011010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011010100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011010100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011011010100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011011010101000) && ({row_reg, col_reg}<16'b0011011010101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011010101011) && ({row_reg, col_reg}<16'b0011011010101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011011010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011010101110) && ({row_reg, col_reg}<16'b0011011010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011010110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011011010110011) && ({row_reg, col_reg}<16'b0011011010110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011011010110110) && ({row_reg, col_reg}<16'b0011011010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011010111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011011010111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011010111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011011010111100) && ({row_reg, col_reg}<16'b0011011010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011011010111110) && ({row_reg, col_reg}<16'b0011011011000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011011000100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0011011011000101) && ({row_reg, col_reg}<16'b0011011011000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011011011000111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011011011001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011011001001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0011011011001010) && ({row_reg, col_reg}<16'b0011011011001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011011011001100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011011011001101)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011011011001110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011011011001111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011011011010000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0011011011010001) && ({row_reg, col_reg}<16'b0011011011010011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011011011010011)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011011011010100)) color_data = 12'b100001110101;
		if(({row_reg, col_reg}==16'b0011011011010101)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011011011010110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011011011010111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011011011011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011011011011001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0011011011011010) && ({row_reg, col_reg}<16'b0011011011011100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011011011011100) && ({row_reg, col_reg}<16'b0011011011011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011011011011110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0011011011011111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011011011100000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011011011100001)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}>=16'b0011011011100010) && ({row_reg, col_reg}<16'b0011011011100100)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==16'b0011011011100100)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011011011100101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0011011011100110) && ({row_reg, col_reg}<16'b0011011011101000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011011011101000) && ({row_reg, col_reg}<16'b0011011011101010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011011011101010)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0011011011101011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011011011101100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011011011101101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011011011101110)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011011011101111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011011011110000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0011011011110001) && ({row_reg, col_reg}<16'b0011011011110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011011011110011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0011011011110100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011011011110101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011011011110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011011011110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011011011111000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011011011111001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011011011111010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011011011111011)) color_data = 12'b100001110101;
		if(({row_reg, col_reg}==16'b0011011011111100)) color_data = 12'b100110000110;
		if(({row_reg, col_reg}==16'b0011011011111101)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==16'b0011011011111110)) color_data = 12'b011001010100;

		if(({row_reg, col_reg}==16'b0011011011111111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011011100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011100000001) && ({row_reg, col_reg}<16'b0011011100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011100000110) && ({row_reg, col_reg}<16'b0011011100001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011011100001001) && ({row_reg, col_reg}<16'b0011011100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011100001100) && ({row_reg, col_reg}<16'b0011011100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011100010010) && ({row_reg, col_reg}<16'b0011011101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011011101100001) && ({row_reg, col_reg}<16'b0011011101100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011101100011) && ({row_reg, col_reg}<16'b0011011101100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011101100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011101100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011101100111) && ({row_reg, col_reg}<16'b0011011101101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011101101001) && ({row_reg, col_reg}<16'b0011011101101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011101101011) && ({row_reg, col_reg}<16'b0011011101101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011101101101) && ({row_reg, col_reg}<16'b0011011101110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011101110101) && ({row_reg, col_reg}<16'b0011011101110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011101110111) && ({row_reg, col_reg}<16'b0011011101111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011101111100) && ({row_reg, col_reg}<16'b0011011101111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011101111110) && ({row_reg, col_reg}<16'b0011011110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011110000001) && ({row_reg, col_reg}<16'b0011011110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011011110010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011110010101) && ({row_reg, col_reg}<16'b0011011110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011011110010111) && ({row_reg, col_reg}<16'b0011011110011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011110011001) && ({row_reg, col_reg}<16'b0011011110011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011011110011100) && ({row_reg, col_reg}<16'b0011011110100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011110100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011011110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011011110100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011011110100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011011110100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011011110101000) && ({row_reg, col_reg}<16'b0011011110101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011011110101011) && ({row_reg, col_reg}<16'b0011011110101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011011110101110) && ({row_reg, col_reg}<16'b0011011110110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011110110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011011110110011) && ({row_reg, col_reg}<16'b0011011110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011011110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011011110110110) && ({row_reg, col_reg}<16'b0011011110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011011110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011011110111001) && ({row_reg, col_reg}<16'b0011011110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011011110111011) && ({row_reg, col_reg}<16'b0011011110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011011110111110) && ({row_reg, col_reg}<16'b0011011111000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011011111000100) && ({row_reg, col_reg}<16'b0011011111001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011011111001000) && ({row_reg, col_reg}<16'b0011011111001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011011111001010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0011011111001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0011011111001100) && ({row_reg, col_reg}<16'b0011011111001110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011011111001110) && ({row_reg, col_reg}<16'b0011011111010000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011011111010000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011011111010001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011011111010010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011011111010011)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}>=16'b0011011111010100) && ({row_reg, col_reg}<16'b0011011111010110)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011011111010110)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011011111010111)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}>=16'b0011011111011000) && ({row_reg, col_reg}<16'b0011011111011011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011011111011011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011011111011100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011011111011101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0011011111011110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011011111011111)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011011111100000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011011111100001)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011011111100010)) color_data = 12'b101111001001;
		if(({row_reg, col_reg}==16'b0011011111100011)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011011111100100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011011111100101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0011011111100110) && ({row_reg, col_reg}<16'b0011011111101011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011011111101011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011011111101100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011011111101101)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011011111101110)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011011111101111)) color_data = 12'b101010111001;
		if(({row_reg, col_reg}==16'b0011011111110000)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011011111110001)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=16'b0011011111110010) && ({row_reg, col_reg}<16'b0011011111110100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011011111110100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011011111110101)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0011011111110110)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0011011111110111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011011111111000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011011111111001)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011011111111010)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011011111111011)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011011111111100)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011011111111101)) color_data = 12'b100110101000;
		if(({row_reg, col_reg}==16'b0011011111111110)) color_data = 12'b011101110110;

		if(({row_reg, col_reg}==16'b0011011111111111)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0011100000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100000000001) && ({row_reg, col_reg}<16'b0011100000000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100000000011) && ({row_reg, col_reg}<16'b0011100000000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011100000000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100000000110) && ({row_reg, col_reg}<16'b0011100000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100000001001) && ({row_reg, col_reg}<16'b0011100000001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100000001101) && ({row_reg, col_reg}<16'b0011100000010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100000010010) && ({row_reg, col_reg}<16'b0011100001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011100001100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100001100010) && ({row_reg, col_reg}<16'b0011100001100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100001100100) && ({row_reg, col_reg}<16'b0011100001100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100001100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100001100111) && ({row_reg, col_reg}<16'b0011100001101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100001101001) && ({row_reg, col_reg}<16'b0011100001101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100001101011) && ({row_reg, col_reg}<16'b0011100001101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100001101101) && ({row_reg, col_reg}<16'b0011100001101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100001101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011100001110000) && ({row_reg, col_reg}<16'b0011100001110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100001110101) && ({row_reg, col_reg}<16'b0011100001110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100001110111) && ({row_reg, col_reg}<16'b0011100001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100001111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100001111101) && ({row_reg, col_reg}<16'b0011100001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011100010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100010000001) && ({row_reg, col_reg}<16'b0011100010010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011100010010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100010010100) && ({row_reg, col_reg}<16'b0011100010010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100010010110) && ({row_reg, col_reg}<16'b0011100010011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100010011000) && ({row_reg, col_reg}<16'b0011100010011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100010011010) && ({row_reg, col_reg}<16'b0011100010011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011100010011100) && ({row_reg, col_reg}<16'b0011100010100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100010100001) && ({row_reg, col_reg}<16'b0011100010100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100010100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011100010100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011100010100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011100010101000) && ({row_reg, col_reg}<16'b0011100010101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100010101011) && ({row_reg, col_reg}<16'b0011100010101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011100010101110) && ({row_reg, col_reg}<16'b0011100010110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100010110011) && ({row_reg, col_reg}<16'b0011100010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011100010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011100010110110) && ({row_reg, col_reg}<16'b0011100010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100010111001) && ({row_reg, col_reg}<16'b0011100010111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011100010111011) && ({row_reg, col_reg}<16'b0011100010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100010111110) && ({row_reg, col_reg}<16'b0011100011000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011100011000111) && ({row_reg, col_reg}<16'b0011100011001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100011001001) && ({row_reg, col_reg}<16'b0011100011001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011100011001011) && ({row_reg, col_reg}<16'b0011100011001110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011100011001110) && ({row_reg, col_reg}<16'b0011100011010001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011100011010001)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011100011010010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011100011010011)) color_data = 12'b100110101000;
		if(({row_reg, col_reg}==16'b0011100011010100)) color_data = 12'b101111001001;
		if(({row_reg, col_reg}==16'b0011100011010101)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==16'b0011100011010110)) color_data = 12'b101010111000;
		if(({row_reg, col_reg}==16'b0011100011010111)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011100011011000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011100011011001)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=16'b0011100011011010) && ({row_reg, col_reg}<16'b0011100011011100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011100011011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011100011011101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011100011011110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011100011011111)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011100011100000)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011100011100001)) color_data = 12'b101111001001;
		if(({row_reg, col_reg}==16'b0011100011100010)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==16'b0011100011100011)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011100011100100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011100011100101)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0011100011100110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011100011100111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0011100011101000) && ({row_reg, col_reg}<16'b0011100011101010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011100011101010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011100011101011)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011100011101100)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=16'b0011100011101101) && ({row_reg, col_reg}<16'b0011100011101111)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==16'b0011100011101111)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011100011110000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011100011110001)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011100011110010)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011100011110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011100011110100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011100011110101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011100011110110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011100011110111)) color_data = 12'b011110000110;
		if(({row_reg, col_reg}>=16'b0011100011111000) && ({row_reg, col_reg}<16'b0011100011111010)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011100011111010)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}>=16'b0011100011111011) && ({row_reg, col_reg}<16'b0011100011111101)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==16'b0011100011111101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011100011111110)) color_data = 12'b010101010011;

		if(({row_reg, col_reg}==16'b0011100011111111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0011100100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100100000001) && ({row_reg, col_reg}<16'b0011100100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100100000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011100100000111) && ({row_reg, col_reg}<16'b0011100100001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100100001001) && ({row_reg, col_reg}<16'b0011100100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100100001011) && ({row_reg, col_reg}<16'b0011100100010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100100010010) && ({row_reg, col_reg}<16'b0011100101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011100101100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100101100010) && ({row_reg, col_reg}<16'b0011100101100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100101100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100101100101) && ({row_reg, col_reg}<16'b0011100101101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100101101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100101101001) && ({row_reg, col_reg}<16'b0011100101110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100101110101) && ({row_reg, col_reg}<16'b0011100101111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100101111000) && ({row_reg, col_reg}<16'b0011100110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011100110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100110000010) && ({row_reg, col_reg}<16'b0011100110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011100110010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011100110010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100110010110) && ({row_reg, col_reg}<16'b0011100110011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100110011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011100110011001) && ({row_reg, col_reg}<16'b0011100110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011100110011101) && ({row_reg, col_reg}<16'b0011100110100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100110100001) && ({row_reg, col_reg}<16'b0011100110100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100110100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011100110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100110100101) && ({row_reg, col_reg}<16'b0011100110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100110101000) && ({row_reg, col_reg}<16'b0011100110101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100110101011) && ({row_reg, col_reg}<16'b0011100110101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011100110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011100110101110) && ({row_reg, col_reg}<16'b0011100110110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011100110110011) && ({row_reg, col_reg}<16'b0011100110110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011100110110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011100110110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011100110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100110111001) && ({row_reg, col_reg}<16'b0011100110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011100110111011) && ({row_reg, col_reg}<16'b0011100110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100110111110) && ({row_reg, col_reg}<16'b0011100111000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011100111000111) && ({row_reg, col_reg}<16'b0011100111001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011100111001001) && ({row_reg, col_reg}<16'b0011100111001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011100111001100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011100111001101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011100111001110)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0011100111001111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0011100111010000) && ({row_reg, col_reg}<16'b0011100111010010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011100111010010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011100111010011)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011100111010100)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==16'b0011100111010101)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011100111010110)) color_data = 12'b110011001001;
		if(({row_reg, col_reg}==16'b0011100111010111)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011100111011000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=16'b0011100111011001) && ({row_reg, col_reg}<16'b0011100111011100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011100111011100)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011100111011101)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0011100111011110)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011100111011111)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011100111100000)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011100111100001)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==16'b0011100111100010)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011100111100011)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011100111100100)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}>=16'b0011100111100101) && ({row_reg, col_reg}<16'b0011100111101001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011100111101001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011100111101010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011100111101011)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==16'b0011100111101100)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011100111101101)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011100111101110)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011100111101111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011100111110000)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011100111110001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0011100111110010) && ({row_reg, col_reg}<16'b0011100111110101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011100111110101)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011100111110110)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==16'b0011100111110111)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011100111111000)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011100111111001)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011100111111010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=16'b0011100111111011) && ({row_reg, col_reg}<16'b0011100111111101)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}>=16'b0011100111111101) && ({row_reg, col_reg}<16'b0011100111111111)) color_data = 12'b010101010100;

		if(({row_reg, col_reg}==16'b0011100111111111)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011101000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011101000000001) && ({row_reg, col_reg}<16'b0011101000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101000000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011101000000111) && ({row_reg, col_reg}<16'b0011101000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101000001001) && ({row_reg, col_reg}<16'b0011101000001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011101000001011) && ({row_reg, col_reg}<16'b0011101000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101000001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011101000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101000010010) && ({row_reg, col_reg}<16'b0011101001100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011101001100010) && ({row_reg, col_reg}<16'b0011101001110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101001110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011101001110100) && ({row_reg, col_reg}<16'b0011101001110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101001110110) && ({row_reg, col_reg}<16'b0011101001111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011101001111000) && ({row_reg, col_reg}<16'b0011101001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101001111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101001111100) && ({row_reg, col_reg}<16'b0011101010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101010000010) && ({row_reg, col_reg}<16'b0011101010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011101010010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101010010101) && ({row_reg, col_reg}<16'b0011101010011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011101010011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101010011001) && ({row_reg, col_reg}<16'b0011101010011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011101010011101) && ({row_reg, col_reg}<16'b0011101010100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101010100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101010100001) && ({row_reg, col_reg}<16'b0011101010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101010100011) && ({row_reg, col_reg}<16'b0011101010100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011101010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101010100110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011101010100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011101010101000) && ({row_reg, col_reg}<16'b0011101010101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011101010101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011101010101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101010101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011101010101101) && ({row_reg, col_reg}<16'b0011101010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011101010110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101010110011) && ({row_reg, col_reg}<16'b0011101010110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101010110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011101010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011101010110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011101010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101010111001) && ({row_reg, col_reg}<16'b0011101010111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011101010111011) && ({row_reg, col_reg}<16'b0011101010111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101010111111) && ({row_reg, col_reg}<16'b0011101011000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101011000011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011101011000100) && ({row_reg, col_reg}<16'b0011101011000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011101011000111) && ({row_reg, col_reg}<16'b0011101011001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101011001001) && ({row_reg, col_reg}<16'b0011101011001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101011001100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011101011001101)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011101011001110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011101011001111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011101011010000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0011101011010001) && ({row_reg, col_reg}<16'b0011101011010011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011101011010011)) color_data = 12'b010101100100;
		if(({row_reg, col_reg}==16'b0011101011010100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011101011010101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==16'b0011101011010110)) color_data = 12'b101111001001;
		if(({row_reg, col_reg}==16'b0011101011010111)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011101011011000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011101011011001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0011101011011010) && ({row_reg, col_reg}<16'b0011101011011100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011101011011100)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011101011011101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011101011011110)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011101011011111)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}>=16'b0011101011100000) && ({row_reg, col_reg}<16'b0011101011100010)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011101011100010)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011101011100011)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}>=16'b0011101011100100) && ({row_reg, col_reg}<16'b0011101011101000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011101011101000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011101011101001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=16'b0011101011101010) && ({row_reg, col_reg}<16'b0011101011101100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011101011101100)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011101011101101)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011101011101110)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=16'b0011101011101111) && ({row_reg, col_reg}<16'b0011101011110001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011101011110001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0011101011110010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011101011110011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011101011110100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011101011110101)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011101011110110)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011101011110111)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011101011111000)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011101011111001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011101011111010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011101011111011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011101011111100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011101011111101)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011101011111110)) color_data = 12'b100010000110;

		if(({row_reg, col_reg}==16'b0011101011111111)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011101100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011101100000001) && ({row_reg, col_reg}<16'b0011101100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101100000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011101100000111) && ({row_reg, col_reg}<16'b0011101100001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101100001001) && ({row_reg, col_reg}<16'b0011101100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011101100001011) && ({row_reg, col_reg}<16'b0011101100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101100001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011101100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101100010001) && ({row_reg, col_reg}<16'b0011101101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011101101100011) && ({row_reg, col_reg}<16'b0011101101101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101101101110) && ({row_reg, col_reg}<16'b0011101101110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101101110100) && ({row_reg, col_reg}<16'b0011101101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101101110110) && ({row_reg, col_reg}<16'b0011101110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101110000010) && ({row_reg, col_reg}<16'b0011101110010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011101110010101) && ({row_reg, col_reg}<16'b0011101110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011101110010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011101110011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011101110011001) && ({row_reg, col_reg}<16'b0011101110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011101110011101) && ({row_reg, col_reg}<16'b0011101110100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101110100000) && ({row_reg, col_reg}<16'b0011101110100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011101110100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011101110100011) && ({row_reg, col_reg}<16'b0011101110100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011101110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011101110100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011101110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011101110101001) && ({row_reg, col_reg}<16'b0011101110101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011101110101011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0011101110101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011101110101101) && ({row_reg, col_reg}<16'b0011101110110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011101110110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101110110011) && ({row_reg, col_reg}<16'b0011101110110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101110110110) && ({row_reg, col_reg}<16'b0011101110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011101110111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011101110111001) && ({row_reg, col_reg}<16'b0011101110111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101110111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011101110111100) && ({row_reg, col_reg}<16'b0011101110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011101110111110) && ({row_reg, col_reg}<16'b0011101111000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101111000011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011101111000100) && ({row_reg, col_reg}<16'b0011101111000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011101111000110) && ({row_reg, col_reg}<16'b0011101111001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101111001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011101111001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011101111001100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011101111001101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011101111001110)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011101111001111)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==16'b0011101111010000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011101111010001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011101111010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011101111010011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011101111010100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011101111010101)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011101111010110)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011101111010111)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011101111011000)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=16'b0011101111011001) && ({row_reg, col_reg}<16'b0011101111011100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011101111011100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011101111011101)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0011101111011110)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011101111011111)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011101111100000)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011101111100001)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011101111100010)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011101111100011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011101111100100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011101111100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011101111100110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011101111100111)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0011101111101000)) color_data = 12'b011110000110;
		if(({row_reg, col_reg}==16'b0011101111101001)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011101111101010)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011101111101011)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011101111101100)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011101111101101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011101111101110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011101111101111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0011101111110000) && ({row_reg, col_reg}<16'b0011101111110010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011101111110010)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}>=16'b0011101111110011) && ({row_reg, col_reg}<16'b0011101111110101)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==16'b0011101111110101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011101111110110)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011101111110111)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011101111111000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0011101111111001) && ({row_reg, col_reg}<16'b0011101111111011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0011101111111011) && ({row_reg, col_reg}<16'b0011101111111101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011101111111101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011101111111110)) color_data = 12'b101110111001;

		if(({row_reg, col_reg}==16'b0011101111111111)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==16'b0011110000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110000000001) && ({row_reg, col_reg}<16'b0011110000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110000000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110000000110) && ({row_reg, col_reg}<16'b0011110000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110000001001) && ({row_reg, col_reg}<16'b0011110000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110000001100) && ({row_reg, col_reg}<16'b0011110000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110000001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011110000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110000010010) && ({row_reg, col_reg}<16'b0011110001100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011110001100100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110001100101) && ({row_reg, col_reg}<16'b0011110001101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110001101010) && ({row_reg, col_reg}<16'b0011110001110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110001110000) && ({row_reg, col_reg}<16'b0011110001110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110001110100) && ({row_reg, col_reg}<16'b0011110001110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110001110110) && ({row_reg, col_reg}<16'b0011110001111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110001111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011110001111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110001111011) && ({row_reg, col_reg}<16'b0011110001111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110001111101) && ({row_reg, col_reg}<16'b0011110010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110010000001) && ({row_reg, col_reg}<16'b0011110010010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011110010010101) && ({row_reg, col_reg}<16'b0011110010011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110010011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110010011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011110010011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011110010011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011110010011100) && ({row_reg, col_reg}<16'b0011110010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110010100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011110010100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011110010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011110010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011110010100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011110010101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110010101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110010101010) && ({row_reg, col_reg}<16'b0011110010101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011110010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110010101110) && ({row_reg, col_reg}<16'b0011110010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110010110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011110010110011) && ({row_reg, col_reg}<16'b0011110010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011110010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011110010110110) && ({row_reg, col_reg}<16'b0011110010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110010111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011110010111001) && ({row_reg, col_reg}<16'b0011110010111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011110010111100) && ({row_reg, col_reg}<16'b0011110010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110010111110) && ({row_reg, col_reg}<16'b0011110011000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110011000011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011110011000100) && ({row_reg, col_reg}<16'b0011110011000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011110011000110) && ({row_reg, col_reg}<16'b0011110011001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011110011001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011110011001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011110011001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110011001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011110011001100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011110011001101)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011110011001110)) color_data = 12'b100010010111;
		if(({row_reg, col_reg}==16'b0011110011001111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011110011010000)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}>=16'b0011110011010001) && ({row_reg, col_reg}<16'b0011110011010100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011110011010100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011110011010101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011110011010110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011110011010111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011110011011000)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==16'b0011110011011001)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011110011011010)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011110011011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0011110011011100) && ({row_reg, col_reg}<16'b0011110011011110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011110011011110)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}>=16'b0011110011011111) && ({row_reg, col_reg}<16'b0011110011100001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011110011100001)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011110011100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011110011100011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011110011100100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011110011100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011110011100110)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0011110011100111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011110011101000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011110011101001)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011110011101010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011110011101011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011110011101100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0011110011101101) && ({row_reg, col_reg}<16'b0011110011101111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011110011101111)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}>=16'b0011110011110000) && ({row_reg, col_reg}<16'b0011110011110010)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011110011110010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011110011110011)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0011110011110100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0011110011110101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011110011110110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011110011110111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011110011111000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011110011111001)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==16'b0011110011111010)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=16'b0011110011111011) && ({row_reg, col_reg}<16'b0011110011111101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011110011111101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==16'b0011110011111110)) color_data = 12'b110011001001;

		if(({row_reg, col_reg}==16'b0011110011111111)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011110100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110100000001) && ({row_reg, col_reg}<16'b0011110100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110100000101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011110100000110) && ({row_reg, col_reg}<16'b0011110100001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011110100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110100001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110100001011) && ({row_reg, col_reg}<16'b0011110100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110100001101) && ({row_reg, col_reg}<16'b0011110100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110100001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011110100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110100010010) && ({row_reg, col_reg}<16'b0011110100110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011110100110001) && ({row_reg, col_reg}<16'b0011110100110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110100110011) && ({row_reg, col_reg}<16'b0011110101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011110101100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110101100100) && ({row_reg, col_reg}<16'b0011110101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110101101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011110101101100) && ({row_reg, col_reg}<16'b0011110101101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110101101110) && ({row_reg, col_reg}<16'b0011110101110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110101110100) && ({row_reg, col_reg}<16'b0011110101110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011110101110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110101111000) && ({row_reg, col_reg}<16'b0011110101111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110101111100) && ({row_reg, col_reg}<16'b0011110101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011110101111110) && ({row_reg, col_reg}<16'b0011110110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110110000010) && ({row_reg, col_reg}<16'b0011110110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011110110010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011110110010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110110010110) && ({row_reg, col_reg}<16'b0011110110011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011110110011000) && ({row_reg, col_reg}<16'b0011110110011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110110011101) && ({row_reg, col_reg}<16'b0011110110011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110110100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011110110100001) && ({row_reg, col_reg}<16'b0011110110100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011110110100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011110110100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011110110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011110110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011110110101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110110101010) && ({row_reg, col_reg}<16'b0011110110101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011110110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110110101110) && ({row_reg, col_reg}<16'b0011110110110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011110110110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011110110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011110110110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110110110110) && ({row_reg, col_reg}<16'b0011110110111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011110110111000) && ({row_reg, col_reg}<16'b0011110110111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011110110111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011110110111100) && ({row_reg, col_reg}<16'b0011110110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110110111110) && ({row_reg, col_reg}<16'b0011110111000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110111000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110111000111) && ({row_reg, col_reg}<16'b0011110111001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011110111001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011110111001010) && ({row_reg, col_reg}<16'b0011110111001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011110111001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0011110111001101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011110111001110)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011110111001111)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0011110111010000)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011110111010001)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011110111010010)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011110111010011)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011110111010100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011110111010101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011110111010110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011110111010111)) color_data = 12'b010101100100;
		if(({row_reg, col_reg}==16'b0011110111011000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011110111011001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0011110111011010) && ({row_reg, col_reg}<16'b0011110111011100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011110111011100)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0011110111011101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011110111011110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011110111011111)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011110111100000)) color_data = 12'b010101100100;
		if(({row_reg, col_reg}==16'b0011110111100001)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011110111100010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011110111100011)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0011110111100100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011110111100101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011110111100110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0011110111100111) && ({row_reg, col_reg}<16'b0011110111101010)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011110111101010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011110111101011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011110111101100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0011110111101101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0011110111101110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011110111101111)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}>=16'b0011110111110000) && ({row_reg, col_reg}<16'b0011110111110010)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011110111110010)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011110111110011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0011110111110100) && ({row_reg, col_reg}<16'b0011110111110110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011110111110110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011110111110111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011110111111000)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011110111111001)) color_data = 12'b101111001001;
		if(({row_reg, col_reg}==16'b0011110111111010)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011110111111011)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011110111111100)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011110111111101)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011110111111110)) color_data = 12'b110011011010;

		if(({row_reg, col_reg}==16'b0011110111111111)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011111000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111000000001) && ({row_reg, col_reg}<16'b0011111000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111000000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011111000000110) && ({row_reg, col_reg}<16'b0011111000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011111000001010) && ({row_reg, col_reg}<16'b0011111000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111000001101) && ({row_reg, col_reg}<16'b0011111000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111000001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011111000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111000010001) && ({row_reg, col_reg}<16'b0011111000011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111000011011) && ({row_reg, col_reg}<16'b0011111000011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111000011111) && ({row_reg, col_reg}<16'b0011111000101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111000101000) && ({row_reg, col_reg}<16'b0011111000101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111000101010) && ({row_reg, col_reg}<16'b0011111000110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011111000110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011111000110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111000110011) && ({row_reg, col_reg}<16'b0011111000110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111000110110) && ({row_reg, col_reg}<16'b0011111000111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111000111000) && ({row_reg, col_reg}<16'b0011111000111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111000111010) && ({row_reg, col_reg}<16'b0011111001001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111001001001) && ({row_reg, col_reg}<16'b0011111001001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111001001101) && ({row_reg, col_reg}<16'b0011111001010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011111001010111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111001011000) && ({row_reg, col_reg}<16'b0011111001011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111001011010) && ({row_reg, col_reg}<16'b0011111001011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111001011100) && ({row_reg, col_reg}<16'b0011111001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011111001100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111001100100) && ({row_reg, col_reg}<16'b0011111001101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111001101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011111001101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111001101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011111001101011)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==16'b0011111001101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111001101101) && ({row_reg, col_reg}<16'b0011111001110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111001110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011111001110010) && ({row_reg, col_reg}<16'b0011111001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111001111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111001111100) && ({row_reg, col_reg}<16'b0011111001111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011111001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111001111111) && ({row_reg, col_reg}<16'b0011111010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111010000010) && ({row_reg, col_reg}<16'b0011111010010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111010010011) && ({row_reg, col_reg}<16'b0011111010010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111010010101) && ({row_reg, col_reg}<16'b0011111010010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111010010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111010011000) && ({row_reg, col_reg}<16'b0011111010011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111010011101) && ({row_reg, col_reg}<16'b0011111010011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011111010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111010100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111010100001) && ({row_reg, col_reg}<16'b0011111010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111010100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011111010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111010100110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011111010100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011111010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011111010101001) && ({row_reg, col_reg}<16'b0011111010101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011111010101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011111010101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011111010101101) && ({row_reg, col_reg}<16'b0011111010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011111010110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011111010110011) && ({row_reg, col_reg}<16'b0011111010110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111010110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011111010110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111010111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011111010111001) && ({row_reg, col_reg}<16'b0011111010111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011111010111011) && ({row_reg, col_reg}<16'b0011111010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011111010111110) && ({row_reg, col_reg}<16'b0011111011000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111011000001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0011111011000010) && ({row_reg, col_reg}<16'b0011111011000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011111011000110) && ({row_reg, col_reg}<16'b0011111011001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011111011001001) && ({row_reg, col_reg}<16'b0011111011001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111011001011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011111011001100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0011111011001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011111011001110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0011111011001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011111011010000)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==16'b0011111011010001)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011111011010010)) color_data = 12'b110111011011;
		if(({row_reg, col_reg}==16'b0011111011010011)) color_data = 12'b101110111000;
		if(({row_reg, col_reg}==16'b0011111011010100)) color_data = 12'b011001110101;
		if(({row_reg, col_reg}>=16'b0011111011010101) && ({row_reg, col_reg}<16'b0011111011010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011111011010111) && ({row_reg, col_reg}<16'b0011111011011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111011011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011111011011011) && ({row_reg, col_reg}<16'b0011111011011110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111011011110)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0011111011011111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011111011100000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111011100001)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}>=16'b0011111011100010) && ({row_reg, col_reg}<16'b0011111011100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011111011100101) && ({row_reg, col_reg}<16'b0011111011101100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011111011101100) && ({row_reg, col_reg}<16'b0011111011101110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111011101110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011111011101111)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0011111011110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0011111011110001) && ({row_reg, col_reg}<16'b0011111011110110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011111011110110)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011111011110111)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011111011111000)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==16'b0011111011111001)) color_data = 12'b110010111001;
		if(({row_reg, col_reg}==16'b0011111011111010)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011111011111011)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011111011111100)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0011111011111101)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011111011111110)) color_data = 12'b101010101000;

		if(({row_reg, col_reg}==16'b0011111011111111)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0011111100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111100000001) && ({row_reg, col_reg}<16'b0011111100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111100000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011111100000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0011111100001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111100001010) && ({row_reg, col_reg}<16'b0011111100001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111100001101) && ({row_reg, col_reg}<16'b0011111100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111100001111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0011111100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111100010001) && ({row_reg, col_reg}<16'b0011111100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011111100010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111100010100) && ({row_reg, col_reg}<16'b0011111100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011111100011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011111100011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111100011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111100011101) && ({row_reg, col_reg}<16'b0011111100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011111100101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011111100101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111100101010) && ({row_reg, col_reg}<16'b0011111100110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111100110000) && ({row_reg, col_reg}<16'b0011111100110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111100110010) && ({row_reg, col_reg}<16'b0011111100110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111100110101) && ({row_reg, col_reg}<16'b0011111100111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111100111010) && ({row_reg, col_reg}<16'b0011111101001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111101001010) && ({row_reg, col_reg}<16'b0011111101001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111101001100) && ({row_reg, col_reg}<16'b0011111101011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011111101011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011111101011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111101011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111101011101) && ({row_reg, col_reg}<16'b0011111101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011111101100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011111101100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111101100101) && ({row_reg, col_reg}<16'b0011111101101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011111101101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011111101101011)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==16'b0011111101101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111101101101) && ({row_reg, col_reg}<16'b0011111101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111101110000) && ({row_reg, col_reg}<16'b0011111101110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011111101110011) && ({row_reg, col_reg}<16'b0011111101111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111101111100) && ({row_reg, col_reg}<16'b0011111101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0011111101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111101111111) && ({row_reg, col_reg}<16'b0011111110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111110000010) && ({row_reg, col_reg}<16'b0011111110010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111110010011) && ({row_reg, col_reg}<16'b0011111110010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0011111110010101) && ({row_reg, col_reg}<16'b0011111110010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111110011000) && ({row_reg, col_reg}<16'b0011111110011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111110011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0011111110011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111110011101) && ({row_reg, col_reg}<16'b0011111110011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111110011111) && ({row_reg, col_reg}<16'b0011111110100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0011111110100001) && ({row_reg, col_reg}<16'b0011111110100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011111110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0011111110100110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0011111110100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011111110101000) && ({row_reg, col_reg}<16'b0011111110101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0011111110101010) && ({row_reg, col_reg}<16'b0011111110110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0011111110110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011111110110011) && ({row_reg, col_reg}<16'b0011111110110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111110110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0011111110110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111110110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0011111110111000) && ({row_reg, col_reg}<16'b0011111110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011111110111011) && ({row_reg, col_reg}<16'b0011111110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011111110111110) && ({row_reg, col_reg}<16'b0011111111000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0011111111000110) && ({row_reg, col_reg}<16'b0011111111001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011111111001000) && ({row_reg, col_reg}<16'b0011111111001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111111001011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011111111001100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0011111111001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011111111001110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0011111111001111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011111111010000)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0011111111010001)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011111111010010)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==16'b0011111111010011)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}==16'b0011111111010100)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0011111111010101)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0011111111010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011111111010111) && ({row_reg, col_reg}<16'b0011111111011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0011111111011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0011111111011010) && ({row_reg, col_reg}<16'b0011111111011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0011111111011100) && ({row_reg, col_reg}<16'b0011111111011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0011111111011110)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0011111111011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011111111100000) && ({row_reg, col_reg}<16'b0011111111100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0011111111100010) && ({row_reg, col_reg}<16'b0011111111100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0011111111100110) && ({row_reg, col_reg}<16'b0011111111101100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0011111111101100) && ({row_reg, col_reg}<16'b0011111111101110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111111101110)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0011111111101111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0011111111110000) && ({row_reg, col_reg}<16'b0011111111110010)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0011111111110010) && ({row_reg, col_reg}<16'b0011111111110100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0011111111110100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011111111110101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0011111111110110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0011111111110111)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011111111111000)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==16'b0011111111111001)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0011111111111010)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==16'b0011111111111011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0011111111111100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0011111111111101)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0011111111111110)) color_data = 12'b011101100101;

		if(({row_reg, col_reg}==16'b0011111111111111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100000000000000) && ({row_reg, col_reg}<16'b0100000000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000000000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100000000000110) && ({row_reg, col_reg}<16'b0100000000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000000001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100000000001010) && ({row_reg, col_reg}<16'b0100000000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000000001111) && ({row_reg, col_reg}<16'b0100000000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100000000010001) && ({row_reg, col_reg}<16'b0100000000010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100000000010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000000010100) && ({row_reg, col_reg}<16'b0100000000011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100000000011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100000000011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000000011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000000011101) && ({row_reg, col_reg}<16'b0100000000101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000000101000) && ({row_reg, col_reg}<16'b0100000000101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000000101010) && ({row_reg, col_reg}<16'b0100000000110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000000110000) && ({row_reg, col_reg}<16'b0100000000110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000000110010) && ({row_reg, col_reg}<16'b0100000000110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000000110110) && ({row_reg, col_reg}<16'b0100000000111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000000111000) && ({row_reg, col_reg}<16'b0100000000111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000000111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000000111011) && ({row_reg, col_reg}<16'b0100000001001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000001001010) && ({row_reg, col_reg}<16'b0100000001001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000001001100) && ({row_reg, col_reg}<16'b0100000001011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100000001011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100000001011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000001011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000001011101) && ({row_reg, col_reg}<16'b0100000001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100000001100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100000001100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000001100101) && ({row_reg, col_reg}<16'b0100000001100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100000001100111) && ({row_reg, col_reg}<16'b0100000001101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000001101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100000001101011)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==16'b0100000001101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000001101101) && ({row_reg, col_reg}<16'b0100000001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000001110000) && ({row_reg, col_reg}<16'b0100000001110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100000001110100) && ({row_reg, col_reg}<16'b0100000001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000001111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100000001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100000001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000001111111) && ({row_reg, col_reg}<16'b0100000010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000010000001) && ({row_reg, col_reg}<16'b0100000010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100000010010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000010010101) && ({row_reg, col_reg}<16'b0100000010010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000010010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100000010011000) && ({row_reg, col_reg}<16'b0100000010011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000010011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100000010011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000010011101) && ({row_reg, col_reg}<16'b0100000010011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100000010011111) && ({row_reg, col_reg}<16'b0100000010100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000010100001) && ({row_reg, col_reg}<16'b0100000010100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100000010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000010100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100000010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100000010101001) && ({row_reg, col_reg}<16'b0100000010110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100000010110001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100000010110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100000010110011) && ({row_reg, col_reg}<16'b0100000010110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000010110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100000010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000010110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100000010111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000010111001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100000010111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100000010111011) && ({row_reg, col_reg}<16'b0100000010111101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0100000010111101) && ({row_reg, col_reg}<16'b0100000011000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100000011000101) && ({row_reg, col_reg}<16'b0100000011001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100000011001001) && ({row_reg, col_reg}<16'b0100000011001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000011001011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0100000011001100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0100000011001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100000011001110)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0100000011001111)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100000011010000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100000011010001)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=16'b0100000011010010) && ({row_reg, col_reg}<16'b0100000011010100)) color_data = 12'b100110010111;
		if(({row_reg, col_reg}==16'b0100000011010100)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0100000011010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100000011010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100000011010111) && ({row_reg, col_reg}<16'b0100000011011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100000011011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100000011011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100000011011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100000011011100) && ({row_reg, col_reg}<16'b0100000011100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000011100000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100000011100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000011100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100000011100011) && ({row_reg, col_reg}<16'b0100000011100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000011100110)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0100000011100111) && ({row_reg, col_reg}<16'b0100000011110100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000011110100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0100000011110101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100000011110110)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=16'b0100000011110111) && ({row_reg, col_reg}<16'b0100000011111001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0100000011111001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100000011111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100000011111011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100000011111100)) color_data = 12'b010001010011;

		if(({row_reg, col_reg}>=16'b0100000011111101) && ({row_reg, col_reg}<16'b0100000100000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0100000100000000) && ({row_reg, col_reg}<16'b0100000100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100000100000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000100000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000100001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000100001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100000100001010) && ({row_reg, col_reg}<16'b0100000100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000100001111) && ({row_reg, col_reg}<16'b0100000100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100000100010001) && ({row_reg, col_reg}<16'b0100000100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100000100011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100000100011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000100011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000100011101) && ({row_reg, col_reg}<16'b0100000100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000100101000) && ({row_reg, col_reg}<16'b0100000100101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000100101010) && ({row_reg, col_reg}<16'b0100000100110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000100110000) && ({row_reg, col_reg}<16'b0100000100110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000100110010) && ({row_reg, col_reg}<16'b0100000100110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000100110110) && ({row_reg, col_reg}<16'b0100000100111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000100111001) && ({row_reg, col_reg}<16'b0100000100111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000100111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000100111100) && ({row_reg, col_reg}<16'b0100000101001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000101001010) && ({row_reg, col_reg}<16'b0100000101001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000101001100) && ({row_reg, col_reg}<16'b0100000101011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100000101011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100000101011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000101011100) && ({row_reg, col_reg}<16'b0100000101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000101100011) && ({row_reg, col_reg}<16'b0100000101100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000101100101) && ({row_reg, col_reg}<16'b0100000101100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100000101100111) && ({row_reg, col_reg}<16'b0100000101101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000101101001) && ({row_reg, col_reg}<16'b0100000101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100000101101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000101101101) && ({row_reg, col_reg}<16'b0100000101110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000101110001) && ({row_reg, col_reg}<16'b0100000101110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100000101110111) && ({row_reg, col_reg}<16'b0100000101111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000101111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000101111110) && ({row_reg, col_reg}<16'b0100000110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100000110000001) && ({row_reg, col_reg}<16'b0100000110010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000110010101) && ({row_reg, col_reg}<16'b0100000110011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100000110011000) && ({row_reg, col_reg}<16'b0100000110011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000110011101) && ({row_reg, col_reg}<16'b0100000110011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100000110011111) && ({row_reg, col_reg}<16'b0100000110100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000110100001) && ({row_reg, col_reg}<16'b0100000110100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100000110100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100000110100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100000110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000110100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100000110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100000110101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100000110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000110101011) && ({row_reg, col_reg}<16'b0100000110101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100000110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100000110101110) && ({row_reg, col_reg}<16'b0100000110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100000110110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100000110110001) && ({row_reg, col_reg}<16'b0100000110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100000110110110) && ({row_reg, col_reg}<16'b0100000110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100000110111000) && ({row_reg, col_reg}<16'b0100000110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100000110111011) && ({row_reg, col_reg}<16'b0100000110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100000110111110) && ({row_reg, col_reg}<16'b0100000111000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100000111000110) && ({row_reg, col_reg}<16'b0100000111001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000111001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000111001011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0100000111001100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0100000111001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100000111001110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100000111001111) && ({row_reg, col_reg}<16'b0100000111010010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100000111010010)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0100000111010011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100000111010100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100000111010101)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0100000111010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100000111010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100000111011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100000111011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100000111011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100000111011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100000111011100) && ({row_reg, col_reg}<16'b0100000111011110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000111011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100000111011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000111100000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100000111100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100000111100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100000111100011) && ({row_reg, col_reg}<16'b0100000111100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100000111100101) && ({row_reg, col_reg}<16'b0100000111100111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100000111100111)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0100000111101000) && ({row_reg, col_reg}<16'b0100000111110100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100000111110100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100000111110101)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100000111110110) && ({row_reg, col_reg}<16'b0100000111111000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100000111111000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100000111111001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100000111111010) && ({row_reg, col_reg}<16'b0100000111111100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100000111111100)) color_data = 12'b010101010011;

		if(({row_reg, col_reg}>=16'b0100000111111101) && ({row_reg, col_reg}<16'b0100001000000000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0100001000000000) && ({row_reg, col_reg}<16'b0100001000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001000000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001000000110) && ({row_reg, col_reg}<16'b0100001000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100001000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100001000001010) && ({row_reg, col_reg}<16'b0100001000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001000001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100001000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001000010001) && ({row_reg, col_reg}<16'b0100001000011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100001000011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001000011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001000011101) && ({row_reg, col_reg}<16'b0100001000110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100001000110000) && ({row_reg, col_reg}<16'b0100001000110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100001000110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001000110011) && ({row_reg, col_reg}<16'b0100001000111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001000111000) && ({row_reg, col_reg}<16'b0100001000111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001000111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001000111011) && ({row_reg, col_reg}<16'b0100001001001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100001001001010) && ({row_reg, col_reg}<16'b0100001001001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001001001100) && ({row_reg, col_reg}<16'b0100001001011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100001001011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100001001011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001001011100) && ({row_reg, col_reg}<16'b0100001001100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100001001100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100001001100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001001100100) && ({row_reg, col_reg}<16'b0100001001100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100001001100110) && ({row_reg, col_reg}<16'b0100001001101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001001101011) && ({row_reg, col_reg}<16'b0100001001101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001001101101) && ({row_reg, col_reg}<16'b0100001001110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001001110010) && ({row_reg, col_reg}<16'b0100001001110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100001001110111) && ({row_reg, col_reg}<16'b0100001001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001001111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100001001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100001001111110) && ({row_reg, col_reg}<16'b0100001010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001010000001) && ({row_reg, col_reg}<16'b0100001010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100001010010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001010010101) && ({row_reg, col_reg}<16'b0100001010011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001010011000) && ({row_reg, col_reg}<16'b0100001010011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001010011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100001010011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001010011101) && ({row_reg, col_reg}<16'b0100001010100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100001010100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001010100001) && ({row_reg, col_reg}<16'b0100001010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001010100011) && ({row_reg, col_reg}<16'b0100001010100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100001010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100001010100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001010100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100001010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100001010101001) && ({row_reg, col_reg}<16'b0100001010101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001010101011) && ({row_reg, col_reg}<16'b0100001010101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100001010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001010101110) && ({row_reg, col_reg}<16'b0100001010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100001010110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100001010110001) && ({row_reg, col_reg}<16'b0100001010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001010110011) && ({row_reg, col_reg}<16'b0100001010110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100001010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100001010110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100001010111000) && ({row_reg, col_reg}<16'b0100001010111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001010111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100001010111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100001010111101) && ({row_reg, col_reg}<16'b0100001010111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001010111111) && ({row_reg, col_reg}<16'b0100001011000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100001011000101) && ({row_reg, col_reg}<16'b0100001011001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100001011001000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0100001011001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100001011001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001011001011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0100001011001100) && ({row_reg, col_reg}<16'b0100001011001110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100001011001110) && ({row_reg, col_reg}<16'b0100001011010000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100001011010000) && ({row_reg, col_reg}<16'b0100001011010011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100001011010011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100001011010100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0100001011010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100001011010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100001011010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100001011011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100001011011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001011011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100001011011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001011011100) && ({row_reg, col_reg}<16'b0100001011011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100001011011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100001011100000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100001011100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100001011100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100001011100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100001011100100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0100001011100101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100001011100110)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100001011100111) && ({row_reg, col_reg}<16'b0100001011110110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100001011110110)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100001011110111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0100001011111000) && ({row_reg, col_reg}<16'b0100001011111110)) color_data = 12'b010001000011;

		if(({row_reg, col_reg}>=16'b0100001011111110) && ({row_reg, col_reg}<16'b0100001100000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100001100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001100000001) && ({row_reg, col_reg}<16'b0100001100000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001100000100) && ({row_reg, col_reg}<16'b0100001100000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001100000110) && ({row_reg, col_reg}<16'b0100001100001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100001100001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100001100001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001100001010) && ({row_reg, col_reg}<16'b0100001100001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001100001101) && ({row_reg, col_reg}<16'b0100001100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001100001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100001100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001100010001) && ({row_reg, col_reg}<16'b0100001100011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100001100011011) && ({row_reg, col_reg}<16'b0100001100011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001100011101) && ({row_reg, col_reg}<16'b0100001100110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100001100110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001100110001) && ({row_reg, col_reg}<16'b0100001100110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001100110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100001100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100001100110101) && ({row_reg, col_reg}<16'b0100001100110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001100110111) && ({row_reg, col_reg}<16'b0100001100111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001100111001) && ({row_reg, col_reg}<16'b0100001100111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001100111011) && ({row_reg, col_reg}<16'b0100001101001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100001101001010) && ({row_reg, col_reg}<16'b0100001101001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001101001100) && ({row_reg, col_reg}<16'b0100001101011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100001101011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100001101011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001101011100) && ({row_reg, col_reg}<16'b0100001101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100001101100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100001101100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001101100100) && ({row_reg, col_reg}<16'b0100001101100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100001101100110) && ({row_reg, col_reg}<16'b0100001101101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001101101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001101101100) && ({row_reg, col_reg}<16'b0100001101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001101101110) && ({row_reg, col_reg}<16'b0100001101110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100001101110111) && ({row_reg, col_reg}<16'b0100001101111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001101111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100001101111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100001101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100001101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001110000001) && ({row_reg, col_reg}<16'b0100001110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100001110010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100001110010101) && ({row_reg, col_reg}<16'b0100001110010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001110011000) && ({row_reg, col_reg}<16'b0100001110011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001110011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100001110011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001110011101) && ({row_reg, col_reg}<16'b0100001110100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001110100000) && ({row_reg, col_reg}<16'b0100001110100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001110100010) && ({row_reg, col_reg}<16'b0100001110100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100001110100101) && ({row_reg, col_reg}<16'b0100001110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100001110101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100001110101001) && ({row_reg, col_reg}<16'b0100001110101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100001110101110) && ({row_reg, col_reg}<16'b0100001110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100001110110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100001110110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100001110110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001110110011) && ({row_reg, col_reg}<16'b0100001110110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001110110110) && ({row_reg, col_reg}<16'b0100001110111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100001110111000) && ({row_reg, col_reg}<16'b0100001110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001110111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001110111100) && ({row_reg, col_reg}<16'b0100001110111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100001110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001110111111) && ({row_reg, col_reg}<16'b0100001111000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100001111000110) && ({row_reg, col_reg}<16'b0100001111001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001111001001) && ({row_reg, col_reg}<16'b0100001111001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100001111001100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100001111001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100001111001110) && ({row_reg, col_reg}<16'b0100001111010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100001111010000) && ({row_reg, col_reg}<16'b0100001111010010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100001111010010)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}>=16'b0100001111010011) && ({row_reg, col_reg}<16'b0100001111010101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100001111010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100001111010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100001111010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100001111011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100001111011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100001111011010) && ({row_reg, col_reg}<16'b0100001111011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100001111011100) && ({row_reg, col_reg}<16'b0100001111011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100001111011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100001111100000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100001111100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100001111100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100001111100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100001111100100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0100001111100101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100001111100110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100001111100111) && ({row_reg, col_reg}<16'b0100001111110101)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100001111110101) && ({row_reg, col_reg}<16'b0100001111111001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100001111111001) && ({row_reg, col_reg}<16'b0100001111111011)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100001111111011)) color_data = 12'b010001000011;

		if(({row_reg, col_reg}>=16'b0100001111111100) && ({row_reg, col_reg}<16'b0100010000000000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100010000000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100010000000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010000000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100010000000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100010000000100) && ({row_reg, col_reg}<16'b0100010000001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100010000001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100010000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010000001010) && ({row_reg, col_reg}<16'b0100010000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010000001101) && ({row_reg, col_reg}<16'b0100010000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010000001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100010000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010000010001) && ({row_reg, col_reg}<16'b0100010000110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010000110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010000110001) && ({row_reg, col_reg}<16'b0100010000110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010000110011) && ({row_reg, col_reg}<16'b0100010000111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010000111100) && ({row_reg, col_reg}<16'b0100010001001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010001001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100010001001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010001001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010001001101) && ({row_reg, col_reg}<16'b0100010001011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010001011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100010001011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010001011100) && ({row_reg, col_reg}<16'b0100010001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100010001100011) && ({row_reg, col_reg}<16'b0100010001100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010001100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100010001100110) && ({row_reg, col_reg}<16'b0100010001101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010001101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100010001101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010001101110) && ({row_reg, col_reg}<16'b0100010001110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100010001110111) && ({row_reg, col_reg}<16'b0100010001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010001111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100010001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100010001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010010000001) && ({row_reg, col_reg}<16'b0100010010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010010010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010010010101) && ({row_reg, col_reg}<16'b0100010010010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010010010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010010011000) && ({row_reg, col_reg}<16'b0100010010011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010010011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100010010011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010010011101) && ({row_reg, col_reg}<16'b0100010010011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010010011111) && ({row_reg, col_reg}<16'b0100010010100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010010100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100010010100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100010010100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100010010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100010010100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100010010100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100010010101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100010010101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010010101010) && ({row_reg, col_reg}<16'b0100010010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100010010110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100010010110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100010010110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100010010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010010110101) && ({row_reg, col_reg}<16'b0100010010111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100010010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010010111001) && ({row_reg, col_reg}<16'b0100010010111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100010010111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100010010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100010010111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100010010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010010111111) && ({row_reg, col_reg}<16'b0100010011000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100010011000111) && ({row_reg, col_reg}<16'b0100010011001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010011001001) && ({row_reg, col_reg}<16'b0100010011001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100010011001100) && ({row_reg, col_reg}<16'b0100010011001111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100010011001111) && ({row_reg, col_reg}<16'b0100010011010010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100010011010010)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0100010011010011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100010011010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100010011010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100010011010110) && ({row_reg, col_reg}<16'b0100010011011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010011011100) && ({row_reg, col_reg}<16'b0100010011011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100010011011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100010011100000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100010011100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100010011100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100010011100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100010011100100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0100010011100101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100010011100110) && ({row_reg, col_reg}<16'b0100010011110110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100010011110110)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0100010011110111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100010011111000) && ({row_reg, col_reg}<16'b0100010011111010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100010011111010)) color_data = 12'b010001010011;

		if(({row_reg, col_reg}>=16'b0100010011111011) && ({row_reg, col_reg}<16'b0100010100000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100010100000000) && ({row_reg, col_reg}<16'b0100010100000010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100010100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010100000011) && ({row_reg, col_reg}<16'b0100010100000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100010100000101) && ({row_reg, col_reg}<16'b0100010100000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010100000111) && ({row_reg, col_reg}<16'b0100010100001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100010100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100010100001010) && ({row_reg, col_reg}<16'b0100010100001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010100001101) && ({row_reg, col_reg}<16'b0100010100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010100001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100010100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010100010010) && ({row_reg, col_reg}<16'b0100010100110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010100110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010100110001) && ({row_reg, col_reg}<16'b0100010100110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010100110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100010100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100010100110101) && ({row_reg, col_reg}<16'b0100010100110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010100110111) && ({row_reg, col_reg}<16'b0100010100111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100010100111011) && ({row_reg, col_reg}<16'b0100010100111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010100111101) && ({row_reg, col_reg}<16'b0100010101001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010101001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100010101001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010101001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010101001101) && ({row_reg, col_reg}<16'b0100010101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010101100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100010101100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010101100101) && ({row_reg, col_reg}<16'b0100010101100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100010101100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010101101000) && ({row_reg, col_reg}<16'b0100010101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100010101101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010101101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010101101101) && ({row_reg, col_reg}<16'b0100010101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010101110000) && ({row_reg, col_reg}<16'b0100010101110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100010101110111) && ({row_reg, col_reg}<16'b0100010101111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010101111100) && ({row_reg, col_reg}<16'b0100010101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100010101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100010110000001) && ({row_reg, col_reg}<16'b0100010110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100010110010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100010110010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010110010110) && ({row_reg, col_reg}<16'b0100010110011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010110011000) && ({row_reg, col_reg}<16'b0100010110011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010110011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100010110011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010110011101) && ({row_reg, col_reg}<16'b0100010110011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100010110011111) && ({row_reg, col_reg}<16'b0100010110100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010110100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100010110100010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100010110100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010110100100) && ({row_reg, col_reg}<16'b0100010110100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100010110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100010110100111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0100010110101000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0100010110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100010110101010) && ({row_reg, col_reg}<16'b0100010110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100010110110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100010110110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100010110110010) && ({row_reg, col_reg}<16'b0100010110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100010110110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100010110110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100010110110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100010110111000) && ({row_reg, col_reg}<16'b0100010110111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010110111011) && ({row_reg, col_reg}<16'b0100010110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100010110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010110111110) && ({row_reg, col_reg}<16'b0100010111001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100010111001100) && ({row_reg, col_reg}<16'b0100010111001110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100010111001110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100010111001111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100010111010000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100010111010001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100010111010010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100010111010011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100010111010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100010111010101) && ({row_reg, col_reg}<16'b0100010111010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100010111010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100010111011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100010111011001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100010111011010) && ({row_reg, col_reg}<16'b0100010111011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100010111011100) && ({row_reg, col_reg}<16'b0100010111011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100010111011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100010111100000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100010111100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100010111100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100010111100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100010111100100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0100010111100101) && ({row_reg, col_reg}<16'b0100010111111011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100010111111011) && ({row_reg, col_reg}<16'b0100010111111101)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100010111111101) && ({row_reg, col_reg}<16'b0100010111111111)) color_data = 12'b010001000011;

		if(({row_reg, col_reg}==16'b0100010111111111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100011000000000) && ({row_reg, col_reg}<16'b0100011000000010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100011000000010) && ({row_reg, col_reg}<16'b0100011000000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100011000000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100011000000110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100011000000111) && ({row_reg, col_reg}<16'b0100011000001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100011000001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011000001010) && ({row_reg, col_reg}<16'b0100011000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011000001101) && ({row_reg, col_reg}<16'b0100011000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011000010010) && ({row_reg, col_reg}<16'b0100011000110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100011000110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100011000110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011000110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011000110011) && ({row_reg, col_reg}<16'b0100011000110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100011000110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011000110110) && ({row_reg, col_reg}<16'b0100011001001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100011001001010) && ({row_reg, col_reg}<16'b0100011001001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011001001100) && ({row_reg, col_reg}<16'b0100011001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100011001100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100011001100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011001100101) && ({row_reg, col_reg}<16'b0100011001100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100011001100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011001101000) && ({row_reg, col_reg}<16'b0100011001101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100011001101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011001101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100011001101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011001101110) && ({row_reg, col_reg}<16'b0100011001110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011001110001) && ({row_reg, col_reg}<16'b0100011001110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100011001110111) && ({row_reg, col_reg}<16'b0100011001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011001111100) && ({row_reg, col_reg}<16'b0100011001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011001111110) && ({row_reg, col_reg}<16'b0100011010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011010000001) && ({row_reg, col_reg}<16'b0100011010010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100011010010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100011010010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011010010101) && ({row_reg, col_reg}<16'b0100011010010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011010010111) && ({row_reg, col_reg}<16'b0100011010011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011010011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100011010011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011010011101) && ({row_reg, col_reg}<16'b0100011010011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100011010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011010100000) && ({row_reg, col_reg}<16'b0100011010100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100011010100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100011010100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011010100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100011010100101) && ({row_reg, col_reg}<16'b0100011010100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011010100111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0100011010101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100011010101001) && ({row_reg, col_reg}<16'b0100011010101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011010101011) && ({row_reg, col_reg}<16'b0100011010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100011010110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100011010110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100011010110010) && ({row_reg, col_reg}<16'b0100011010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100011010110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100011010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011010110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100011010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100011010111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100011010111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100011010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100011010111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100011010111110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100011010111111) && ({row_reg, col_reg}<16'b0100011011000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100011011000010) && ({row_reg, col_reg}<16'b0100011011001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011011001011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0100011011001100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100011011001101) && ({row_reg, col_reg}<16'b0100011011010000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100011011010000) && ({row_reg, col_reg}<16'b0100011011010010)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100011011010010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100011011010011) && ({row_reg, col_reg}<16'b0100011011010101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100011011010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100011011010110) && ({row_reg, col_reg}<16'b0100011011011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011011011000) && ({row_reg, col_reg}<16'b0100011011011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100011011011010) && ({row_reg, col_reg}<16'b0100011011011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011011011100) && ({row_reg, col_reg}<16'b0100011011011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011011011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100011011100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011011100001) && ({row_reg, col_reg}<16'b0100011011100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100011011100011) && ({row_reg, col_reg}<16'b0100011011100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100011011100101) && ({row_reg, col_reg}<16'b0100011011110111)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0100011011110111) && ({row_reg, col_reg}<16'b0100011011111001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100011011111001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100011011111010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100011011111011)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100011011111100) && ({row_reg, col_reg}<16'b0100011011111110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100011011111110)) color_data = 12'b001101000010;

		if(({row_reg, col_reg}==16'b0100011011111111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100011100000000) && ({row_reg, col_reg}<16'b0100011100000101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100011100000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011100000110) && ({row_reg, col_reg}<16'b0100011100001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100011100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011100001010) && ({row_reg, col_reg}<16'b0100011100001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011100001101) && ({row_reg, col_reg}<16'b0100011100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100011100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011100010001) && ({row_reg, col_reg}<16'b0100011100110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100011100110000) && ({row_reg, col_reg}<16'b0100011100110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011100110011) && ({row_reg, col_reg}<16'b0100011100110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100011100110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011100110110) && ({row_reg, col_reg}<16'b0100011101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100011101100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100011101100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011101100101) && ({row_reg, col_reg}<16'b0100011101100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100011101100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011101101000) && ({row_reg, col_reg}<16'b0100011101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100011101101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011101101101) && ({row_reg, col_reg}<16'b0100011101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011101110000) && ({row_reg, col_reg}<16'b0100011101110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100011101110101) && ({row_reg, col_reg}<16'b0100011101111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011101111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100011101111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100011101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100011101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100011110000001) && ({row_reg, col_reg}<16'b0100011110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100011110010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011110010101) && ({row_reg, col_reg}<16'b0100011110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011110010111) && ({row_reg, col_reg}<16'b0100011110011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011110011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100011110011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100011110011101) && ({row_reg, col_reg}<16'b0100011110011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100011110011111) && ({row_reg, col_reg}<16'b0100011110100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011110100001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100011110100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100011110100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100011110100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011110100101) && ({row_reg, col_reg}<16'b0100011110101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100011110101001) && ({row_reg, col_reg}<16'b0100011110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100011110101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100011110101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100011110101101) && ({row_reg, col_reg}<16'b0100011110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100011110110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100011110110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100011110110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011110110011) && ({row_reg, col_reg}<16'b0100011110110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100011110110101) && ({row_reg, col_reg}<16'b0100011110111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100011110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011110111001) && ({row_reg, col_reg}<16'b0100011110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011110111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100011110111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100011110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100011110111110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100011110111111) && ({row_reg, col_reg}<16'b0100011111000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100011111000010) && ({row_reg, col_reg}<16'b0100011111001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100011111001011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0100011111001100) && ({row_reg, col_reg}<16'b0100011111001110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100011111001110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100011111001111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100011111010000) && ({row_reg, col_reg}<16'b0100011111010101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100011111010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011111010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011111010111) && ({row_reg, col_reg}<16'b0100011111011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100011111011010) && ({row_reg, col_reg}<16'b0100011111011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100011111011100) && ({row_reg, col_reg}<16'b0100011111011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011111011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100011111100000) && ({row_reg, col_reg}<16'b0100011111100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100011111100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100011111100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011111100100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0100011111100101) && ({row_reg, col_reg}<16'b0100011111111000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100011111111000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100011111111001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100011111111010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100011111111011)) color_data = 12'b010001010011;

		if(({row_reg, col_reg}>=16'b0100011111111100) && ({row_reg, col_reg}<16'b0100100000000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100100000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100000000001) && ({row_reg, col_reg}<16'b0100100000000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100000000100) && ({row_reg, col_reg}<16'b0100100000000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100100000000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100000000111) && ({row_reg, col_reg}<16'b0100100000001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100100000001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100000001010) && ({row_reg, col_reg}<16'b0100100000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100000001110) && ({row_reg, col_reg}<16'b0100100000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100000010001) && ({row_reg, col_reg}<16'b0100100000110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100100000110010) && ({row_reg, col_reg}<16'b0100100000110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100100000110110) && ({row_reg, col_reg}<16'b0100100001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100100001100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100100001100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100001100101) && ({row_reg, col_reg}<16'b0100100001100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100100001100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100001101000) && ({row_reg, col_reg}<16'b0100100001101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100001101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100100001101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100001101110) && ({row_reg, col_reg}<16'b0100100001110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100100001110101) && ({row_reg, col_reg}<16'b0100100001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100001111100) && ({row_reg, col_reg}<16'b0100100001111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100100001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100100001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100100010000001) && ({row_reg, col_reg}<16'b0100100010010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100100010010101) && ({row_reg, col_reg}<16'b0100100010010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100010010111) && ({row_reg, col_reg}<16'b0100100010011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100010011101) && ({row_reg, col_reg}<16'b0100100010011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100010011111) && ({row_reg, col_reg}<16'b0100100010100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100010100001) && ({row_reg, col_reg}<16'b0100100010100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100010100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100100010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100100010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100010100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100100010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100100010101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100010101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100010101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100100010101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100100010101101) && ({row_reg, col_reg}<16'b0100100010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100010110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100100010110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100100010110010) && ({row_reg, col_reg}<16'b0100100010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100100010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100100010110110) && ({row_reg, col_reg}<16'b0100100010111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100100010111000) && ({row_reg, col_reg}<16'b0100100010111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100100010111011) && ({row_reg, col_reg}<16'b0100100010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100010111110) && ({row_reg, col_reg}<16'b0100100011000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100100011000000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0100100011000001) && ({row_reg, col_reg}<16'b0100100011000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100100011000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100011000111) && ({row_reg, col_reg}<16'b0100100011001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100100011001011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0100100011001100) && ({row_reg, col_reg}<16'b0100100011001110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100100011001110)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0100100011001111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100100011010000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100100011010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100100011010010) && ({row_reg, col_reg}<16'b0100100011010101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100100011010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100011010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100011010111) && ({row_reg, col_reg}<16'b0100100011011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100011011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100100011011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100011011100) && ({row_reg, col_reg}<16'b0100100011011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100011011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100100011100000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100100011100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100100011100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100100011100011) && ({row_reg, col_reg}<16'b0100100011111000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100011111000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100100011111001)) color_data = 12'b010101010100;

		if(({row_reg, col_reg}>=16'b0100100011111010) && ({row_reg, col_reg}<16'b0100100100000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100100100000000) && ({row_reg, col_reg}<16'b0100100100000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100100000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100100000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100100000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100100100000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100100000111) && ({row_reg, col_reg}<16'b0100100100001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100100100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100100001010) && ({row_reg, col_reg}<16'b0100100100001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100100001110) && ({row_reg, col_reg}<16'b0100100100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100100010001) && ({row_reg, col_reg}<16'b0100100101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100100101100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100100101100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100101100101) && ({row_reg, col_reg}<16'b0100100101100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100100101100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100101101000) && ({row_reg, col_reg}<16'b0100100101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100101101011) && ({row_reg, col_reg}<16'b0100100101101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100100101101101) && ({row_reg, col_reg}<16'b0100100101110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100101110001) && ({row_reg, col_reg}<16'b0100100101110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100100101110101) && ({row_reg, col_reg}<16'b0100100101111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100100101111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100100101111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100100101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100100101111111) && ({row_reg, col_reg}<16'b0100100110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100110000001) && ({row_reg, col_reg}<16'b0100100110010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100100110010101) && ({row_reg, col_reg}<16'b0100100110011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100110011000) && ({row_reg, col_reg}<16'b0100100110011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100110011101) && ({row_reg, col_reg}<16'b0100100110011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100110100000) && ({row_reg, col_reg}<16'b0100100110100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100100110100010) && ({row_reg, col_reg}<16'b0100100110100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100110100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100100110100110) && ({row_reg, col_reg}<16'b0100100110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100110101000) && ({row_reg, col_reg}<16'b0100100110101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100100110101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100100110101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100100110101101) && ({row_reg, col_reg}<16'b0100100110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100100110110000) && ({row_reg, col_reg}<16'b0100100110110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100100110110011) && ({row_reg, col_reg}<16'b0100100110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100110110101) && ({row_reg, col_reg}<16'b0100100110111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100100110111000) && ({row_reg, col_reg}<16'b0100100110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100100110111011) && ({row_reg, col_reg}<16'b0100100110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100110111110) && ({row_reg, col_reg}<16'b0100100111000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100100111000101) && ({row_reg, col_reg}<16'b0100100111000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100111000111) && ({row_reg, col_reg}<16'b0100100111001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100100111001011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0100100111001100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0100100111001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100100111001110)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0100100111001111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100100111010000) && ({row_reg, col_reg}<16'b0100100111010101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100100111010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100111010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100100111010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100100111011000) && ({row_reg, col_reg}<16'b0100100111011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100100111011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100100111011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100100111011100) && ({row_reg, col_reg}<16'b0100100111011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100111011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100100111100000) && ({row_reg, col_reg}<16'b0100100111100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100100111100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100100111100011) && ({row_reg, col_reg}<16'b0100100111100101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100111100101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0100100111100110) && ({row_reg, col_reg}<16'b0100100111101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100100111101011) && ({row_reg, col_reg}<16'b0100100111101101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0100100111101101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0100100111101110)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0100100111101111) && ({row_reg, col_reg}<16'b0100100111110010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100100111110010) && ({row_reg, col_reg}<16'b0100100111110100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0100100111110100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0100100111110101)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0100100111110110) && ({row_reg, col_reg}<16'b0100100111111000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100100111111000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100100111111001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100100111111010) && ({row_reg, col_reg}<16'b0100100111111101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100100111111101) && ({row_reg, col_reg}<16'b0100100111111111)) color_data = 12'b010001010011;

		if(({row_reg, col_reg}==16'b0100100111111111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100101000000000) && ({row_reg, col_reg}<16'b0100101000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101000000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100101000000111) && ({row_reg, col_reg}<16'b0100101000001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100101000001001) && ({row_reg, col_reg}<16'b0100101000001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101000001011) && ({row_reg, col_reg}<16'b0100101000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101000001111) && ({row_reg, col_reg}<16'b0100101000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101000010001) && ({row_reg, col_reg}<16'b0100101000111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101000111010) && ({row_reg, col_reg}<16'b0100101000111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101000111101) && ({row_reg, col_reg}<16'b0100101001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100101001100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101001100100) && ({row_reg, col_reg}<16'b0100101001100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101001100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100101001100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101001101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101001101001) && ({row_reg, col_reg}<16'b0100101001101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101001101011) && ({row_reg, col_reg}<16'b0100101001101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101001101101) && ({row_reg, col_reg}<16'b0100101001110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101001110001) && ({row_reg, col_reg}<16'b0100101001110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100101001110111) && ({row_reg, col_reg}<16'b0100101001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101001111100) && ({row_reg, col_reg}<16'b0100101001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100101001111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101001111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100101010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101010000010) && ({row_reg, col_reg}<16'b0100101010010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101010010101) && ({row_reg, col_reg}<16'b0100101010011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101010011000) && ({row_reg, col_reg}<16'b0100101010011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101010011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100101010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101010100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100101010100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101010100010) && ({row_reg, col_reg}<16'b0100101010100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100101010100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100101010100110) && ({row_reg, col_reg}<16'b0100101010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101010101000) && ({row_reg, col_reg}<16'b0100101010101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100101010101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100101010101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100101010101101) && ({row_reg, col_reg}<16'b0100101010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101010110000) && ({row_reg, col_reg}<16'b0100101010110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100101010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101010110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101010110110) && ({row_reg, col_reg}<16'b0100101010111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100101010111000) && ({row_reg, col_reg}<16'b0100101010111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100101010111011) && ({row_reg, col_reg}<16'b0100101010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101010111110) && ({row_reg, col_reg}<16'b0100101011000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100101011000110) && ({row_reg, col_reg}<16'b0100101011001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101011001001) && ({row_reg, col_reg}<16'b0100101011001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101011001011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100101011001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0100101011001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100101011001110)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0100101011001111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100101011010000) && ({row_reg, col_reg}<16'b0100101011010010)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100101011010010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100101011010011) && ({row_reg, col_reg}<16'b0100101011010101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100101011010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100101011010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100101011010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100101011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100101011011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101011011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100101011011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101011011100) && ({row_reg, col_reg}<16'b0100101011011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100101011011111) && ({row_reg, col_reg}<16'b0100101011100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100101011100011) && ({row_reg, col_reg}<16'b0100101011101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100101011101000) && ({row_reg, col_reg}<16'b0100101011101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100101011101010) && ({row_reg, col_reg}<16'b0100101011110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100101011110000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100101011110001) && ({row_reg, col_reg}<16'b0100101011111000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100101011111000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100101011111001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100101011111010)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100101011111011) && ({row_reg, col_reg}<16'b0100101011111101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0100101011111101)) color_data = 12'b010001010011;

		if(({row_reg, col_reg}>=16'b0100101011111110) && ({row_reg, col_reg}<16'b0100101100000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100101100000000) && ({row_reg, col_reg}<16'b0100101100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101100000110) && ({row_reg, col_reg}<16'b0100101100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101100001010) && ({row_reg, col_reg}<16'b0100101100001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101100001101) && ({row_reg, col_reg}<16'b0100101100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101100001111) && ({row_reg, col_reg}<16'b0100101100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101100010001) && ({row_reg, col_reg}<16'b0100101100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100101100010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101100010100) && ({row_reg, col_reg}<16'b0100101100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101100111001) && ({row_reg, col_reg}<16'b0100101100111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101100111101) && ({row_reg, col_reg}<16'b0100101101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100101101100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101101100100) && ({row_reg, col_reg}<16'b0100101101101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101101101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101101101001) && ({row_reg, col_reg}<16'b0100101101101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101101101011) && ({row_reg, col_reg}<16'b0100101101101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101101101101) && ({row_reg, col_reg}<16'b0100101101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101101110000) && ({row_reg, col_reg}<16'b0100101101110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100101101110111) && ({row_reg, col_reg}<16'b0100101101111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101101111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100101101111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101101111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100101110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100101110000010) && ({row_reg, col_reg}<16'b0100101110010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101110010101) && ({row_reg, col_reg}<16'b0100101110011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101110011001) && ({row_reg, col_reg}<16'b0100101110011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101110011101) && ({row_reg, col_reg}<16'b0100101110011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101110011111) && ({row_reg, col_reg}<16'b0100101110100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100101110100001) && ({row_reg, col_reg}<16'b0100101110100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100101110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101110100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100101110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101110101000) && ({row_reg, col_reg}<16'b0100101110101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100101110101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101110101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100101110101100) && ({row_reg, col_reg}<16'b0100101110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100101110110000) && ({row_reg, col_reg}<16'b0100101110110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100101110110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101110110011) && ({row_reg, col_reg}<16'b0100101110110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101110110110) && ({row_reg, col_reg}<16'b0100101110111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100101110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101110111001) && ({row_reg, col_reg}<16'b0100101110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100101110111011) && ({row_reg, col_reg}<16'b0100101110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101110111110) && ({row_reg, col_reg}<16'b0100101111000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100101111000110) && ({row_reg, col_reg}<16'b0100101111001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101111001001) && ({row_reg, col_reg}<16'b0100101111001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101111001011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0100101111001100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0100101111001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100101111001110)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100101111001111) && ({row_reg, col_reg}<16'b0100101111010001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100101111010001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100101111010010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100101111010011) && ({row_reg, col_reg}<16'b0100101111010101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100101111010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100101111010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101111010111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==16'b0100101111011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100101111011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100101111011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100101111011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101111011100) && ({row_reg, col_reg}<16'b0100101111011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100101111011111) && ({row_reg, col_reg}<16'b0100101111100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100101111100010) && ({row_reg, col_reg}<16'b0100101111100100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100101111100100) && ({row_reg, col_reg}<16'b0100101111100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100101111100111) && ({row_reg, col_reg}<16'b0100101111101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101111101010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100101111101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100101111101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100101111101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101111101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100101111101111) && ({row_reg, col_reg}<16'b0100101111110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101111110001) && ({row_reg, col_reg}<16'b0100101111110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100101111110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100101111110100) && ({row_reg, col_reg}<16'b0100101111110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100101111110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100101111110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100101111111000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100101111111001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100101111111010)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0100101111111011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0100101111111100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0100101111111101)) color_data = 12'b010101010100;

		if(({row_reg, col_reg}>=16'b0100101111111110) && ({row_reg, col_reg}<16'b0100110000000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100110000000000) && ({row_reg, col_reg}<16'b0100110000000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110000000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100110000000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110000000101) && ({row_reg, col_reg}<16'b0100110000001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100110000001001) && ({row_reg, col_reg}<16'b0100110000001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100110000001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100110000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100110000001101) && ({row_reg, col_reg}<16'b0100110000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110000001111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100110000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110000010001) && ({row_reg, col_reg}<16'b0100110000010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100110000010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110000010100) && ({row_reg, col_reg}<16'b0100110000111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110000111000) && ({row_reg, col_reg}<16'b0100110000111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110000111101) && ({row_reg, col_reg}<16'b0100110001001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110001001011) && ({row_reg, col_reg}<16'b0100110001001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110001001101) && ({row_reg, col_reg}<16'b0100110001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110001100011) && ({row_reg, col_reg}<16'b0100110001101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110001101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100110001101001) && ({row_reg, col_reg}<16'b0100110001101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110001101011) && ({row_reg, col_reg}<16'b0100110001101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100110001101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100110001101110) && ({row_reg, col_reg}<16'b0100110001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110001110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100110001110001) && ({row_reg, col_reg}<16'b0100110001110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110001110101) && ({row_reg, col_reg}<16'b0100110001110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100110001110111) && ({row_reg, col_reg}<16'b0100110001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110001111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110010000010) && ({row_reg, col_reg}<16'b0100110010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100110010010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100110010010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110010010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110010010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110010011000) && ({row_reg, col_reg}<16'b0100110010011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100110010011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110010011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100110010011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110010011101) && ({row_reg, col_reg}<16'b0100110010011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100110010011111) && ({row_reg, col_reg}<16'b0100110010100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110010100010) && ({row_reg, col_reg}<16'b0100110010100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110010100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100110010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100110010100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100110010101000) && ({row_reg, col_reg}<16'b0100110010101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100110010101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110010101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100110010101101) && ({row_reg, col_reg}<16'b0100110010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100110010110000) && ({row_reg, col_reg}<16'b0100110010110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100110010110010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0100110010110011) && ({row_reg, col_reg}<16'b0100110010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100110010110110) && ({row_reg, col_reg}<16'b0100110010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100110010111001) && ({row_reg, col_reg}<16'b0100110010111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100110010111011) && ({row_reg, col_reg}<16'b0100110010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100110010111110) && ({row_reg, col_reg}<16'b0100110011000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100110011000110) && ({row_reg, col_reg}<16'b0100110011001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100110011001001) && ({row_reg, col_reg}<16'b0100110011001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100110011001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100110011001100) && ({row_reg, col_reg}<16'b0100110011001110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100110011001110)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}>=16'b0100110011001111) && ({row_reg, col_reg}<16'b0100110011010001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0100110011010001) && ({row_reg, col_reg}<16'b0100110011010101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100110011010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100110011010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110011010111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==16'b0100110011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100110011011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110011011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100110011011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100110011011100) && ({row_reg, col_reg}<16'b0100110011011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100110011011111) && ({row_reg, col_reg}<16'b0100110011100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100110011100010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100110011100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100110011100100) && ({row_reg, col_reg}<16'b0100110011101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100110011101000) && ({row_reg, col_reg}<16'b0100110011101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100110011101010) && ({row_reg, col_reg}<16'b0100110011101100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100110011101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100110011101101) && ({row_reg, col_reg}<16'b0100110011110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100110011110000) && ({row_reg, col_reg}<16'b0100110011110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100110011110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100110011110100) && ({row_reg, col_reg}<16'b0100110011110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110011110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100110011110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100110011111000) && ({row_reg, col_reg}<16'b0100110011111011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100110011111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0100110011111100) && ({row_reg, col_reg}<16'b0100110011111110)) color_data = 12'b010101010011;

		if(({row_reg, col_reg}>=16'b0100110011111110) && ({row_reg, col_reg}<16'b0100110100000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100110100000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100110100000001) && ({row_reg, col_reg}<16'b0100110100000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110100000011) && ({row_reg, col_reg}<16'b0100110100000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110100000101) && ({row_reg, col_reg}<16'b0100110100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100110100001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100110100001001) && ({row_reg, col_reg}<16'b0100110100001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100110100001011) && ({row_reg, col_reg}<16'b0100110100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100110100001101) && ({row_reg, col_reg}<16'b0100110100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110100010010) && ({row_reg, col_reg}<16'b0100110100110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110100110001) && ({row_reg, col_reg}<16'b0100110100110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110100110011) && ({row_reg, col_reg}<16'b0100110100111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110100111000) && ({row_reg, col_reg}<16'b0100110100111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110100111101) && ({row_reg, col_reg}<16'b0100110101001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110101001011) && ({row_reg, col_reg}<16'b0100110101001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110101001101) && ({row_reg, col_reg}<16'b0100110101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100110101100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100110101100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110101100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100110101100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110101100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100110101100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110101101000) && ({row_reg, col_reg}<16'b0100110101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110101101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110101101100) && ({row_reg, col_reg}<16'b0100110101110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110101110101) && ({row_reg, col_reg}<16'b0100110101110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100110101110111) && ({row_reg, col_reg}<16'b0100110101111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110101111110) && ({row_reg, col_reg}<16'b0100110110000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110110000001) && ({row_reg, col_reg}<16'b0100110110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100110110010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110110010101) && ({row_reg, col_reg}<16'b0100110110011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110110011000) && ({row_reg, col_reg}<16'b0100110110011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110110011011) && ({row_reg, col_reg}<16'b0100110110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110110011101) && ({row_reg, col_reg}<16'b0100110110011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110110100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100110110100001) && ({row_reg, col_reg}<16'b0100110110100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100110110100011) && ({row_reg, col_reg}<16'b0100110110100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100110110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100110110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100110110100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100110110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100110110101001) && ({row_reg, col_reg}<16'b0100110110101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100110110101011) && ({row_reg, col_reg}<16'b0100110110101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100110110101101) && ({row_reg, col_reg}<16'b0100110110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100110110110000) && ({row_reg, col_reg}<16'b0100110110110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100110110110010) && ({row_reg, col_reg}<16'b0100110110110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100110110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100110110110110) && ({row_reg, col_reg}<16'b0100110110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110110111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100110110111001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100110110111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100110110111011) && ({row_reg, col_reg}<16'b0100110110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100110110111110) && ({row_reg, col_reg}<16'b0100110111000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100110111000110) && ({row_reg, col_reg}<16'b0100110111001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100110111001001) && ({row_reg, col_reg}<16'b0100110111001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100110111001011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0100110111001100) && ({row_reg, col_reg}<16'b0100110111001110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0100110111001110)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0100110111001111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100110111010000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100110111010001) && ({row_reg, col_reg}<16'b0100110111010011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100110111010011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100110111010100)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==16'b0100110111010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100110111010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100110111010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100110111011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100110111011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100110111011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100110111011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100110111011100) && ({row_reg, col_reg}<16'b0100110111011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100110111011111) && ({row_reg, col_reg}<16'b0100110111100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100110111100011) && ({row_reg, col_reg}<16'b0100110111101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100110111101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100110111101001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100110111101010) && ({row_reg, col_reg}<16'b0100110111101110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100110111101110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100110111101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100110111110000) && ({row_reg, col_reg}<16'b0100110111111000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100110111111000)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}>=16'b0100110111111001) && ({row_reg, col_reg}<16'b0100110111111100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100110111111100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0100110111111101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100110111111110)) color_data = 12'b010001010011;

		if(({row_reg, col_reg}==16'b0100110111111111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100111000000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100111000000001) && ({row_reg, col_reg}<16'b0100111000000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111000000011) && ({row_reg, col_reg}<16'b0100111000000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111000000101) && ({row_reg, col_reg}<16'b0100111000000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111000000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100111000001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100111000001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100111000001011) && ({row_reg, col_reg}<16'b0100111000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111000010010) && ({row_reg, col_reg}<16'b0100111000111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111000111000) && ({row_reg, col_reg}<16'b0100111000111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111000111101) && ({row_reg, col_reg}<16'b0100111001100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100111001100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100111001100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111001100100) && ({row_reg, col_reg}<16'b0100111001100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100111001100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111001101000) && ({row_reg, col_reg}<16'b0100111001101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111001101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111001101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111001101100) && ({row_reg, col_reg}<16'b0100111001110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111001110010) && ({row_reg, col_reg}<16'b0100111001110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111001110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111001110101) && ({row_reg, col_reg}<16'b0100111001110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100111001110111) && ({row_reg, col_reg}<16'b0100111001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111001111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111001111110) && ({row_reg, col_reg}<16'b0100111010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111010000001) && ({row_reg, col_reg}<16'b0100111010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111010010100) && ({row_reg, col_reg}<16'b0100111010011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111010011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111010011001) && ({row_reg, col_reg}<16'b0100111010011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111010011101) && ({row_reg, col_reg}<16'b0100111010011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100111010011111) && ({row_reg, col_reg}<16'b0100111010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111010100011) && ({row_reg, col_reg}<16'b0100111010100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100111010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100111010100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100111010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100111010101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111010101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100111010101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100111010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111010101110) && ({row_reg, col_reg}<16'b0100111010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100111010110000) && ({row_reg, col_reg}<16'b0100111010110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100111010110011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0100111010110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100111010110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100111010110110) && ({row_reg, col_reg}<16'b0100111010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111010111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100111010111001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0100111010111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100111010111011) && ({row_reg, col_reg}<16'b0100111010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100111010111110) && ({row_reg, col_reg}<16'b0100111011000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100111011000010) && ({row_reg, col_reg}<16'b0100111011000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111011000110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0100111011000111) && ({row_reg, col_reg}<16'b0100111011001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111011001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100111011001011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0100111011001100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0100111011001101) && ({row_reg, col_reg}<16'b0100111011010011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100111011010011) && ({row_reg, col_reg}<16'b0100111011010101)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0100111011010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100111011010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100111011010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100111011011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111011011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100111011011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100111011011100) && ({row_reg, col_reg}<16'b0100111011011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100111011011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100111011100000) && ({row_reg, col_reg}<16'b0100111011100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111011100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0100111011100011) && ({row_reg, col_reg}<16'b0100111011101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100111011101011)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0100111011101100) && ({row_reg, col_reg}<16'b0100111011111000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100111011111000) && ({row_reg, col_reg}<16'b0100111011111010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0100111011111010) && ({row_reg, col_reg}<16'b0100111011111100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100111011111100) && ({row_reg, col_reg}<16'b0100111011111110)) color_data = 12'b010001000011;

		if(({row_reg, col_reg}>=16'b0100111011111110) && ({row_reg, col_reg}<16'b0100111100000000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0100111100000000) && ({row_reg, col_reg}<16'b0100111100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111100000101) && ({row_reg, col_reg}<16'b0100111100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100111100001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100111100001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100111100001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111100001110) && ({row_reg, col_reg}<16'b0100111100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100111100010001) && ({row_reg, col_reg}<16'b0100111100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111100111001) && ({row_reg, col_reg}<16'b0100111100111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111100111101) && ({row_reg, col_reg}<16'b0100111101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0100111101100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100111101100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111101100100) && ({row_reg, col_reg}<16'b0100111101100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100111101100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111101101000) && ({row_reg, col_reg}<16'b0100111101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111101101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111101101100) && ({row_reg, col_reg}<16'b0100111101110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111101110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100111101110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111101110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111101110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111101110101) && ({row_reg, col_reg}<16'b0100111101110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0100111101110111) && ({row_reg, col_reg}<16'b0100111101111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111101111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111101111100) && ({row_reg, col_reg}<16'b0100111101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100111101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0100111110000001) && ({row_reg, col_reg}<16'b0100111110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111110010100) && ({row_reg, col_reg}<16'b0100111110010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100111110010110) && ({row_reg, col_reg}<16'b0100111110011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111110011000) && ({row_reg, col_reg}<16'b0100111110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111110011101) && ({row_reg, col_reg}<16'b0100111110011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100111110011111) && ({row_reg, col_reg}<16'b0100111110100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111110100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0100111110100010) && ({row_reg, col_reg}<16'b0100111110100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100111110100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100111110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100111110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100111110101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111110101011) && ({row_reg, col_reg}<16'b0100111110101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100111110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0100111110101110) && ({row_reg, col_reg}<16'b0100111110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111110110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0100111110110001) && ({row_reg, col_reg}<16'b0100111110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111110110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100111110110101) && ({row_reg, col_reg}<16'b0100111110110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100111110110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100111110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100111110111001) && ({row_reg, col_reg}<16'b0100111110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100111110111011) && ({row_reg, col_reg}<16'b0100111110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100111110111110) && ({row_reg, col_reg}<16'b0100111111000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0100111111000010) && ({row_reg, col_reg}<16'b0100111111000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100111111000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100111111000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100111111000110) && ({row_reg, col_reg}<16'b0100111111001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0100111111001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100111111001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111111001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0100111111001011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0100111111001100) && ({row_reg, col_reg}<16'b0100111111001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0100111111001110) && ({row_reg, col_reg}<16'b0100111111010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100111111010000) && ({row_reg, col_reg}<16'b0100111111010010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100111111010010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100111111010011) && ({row_reg, col_reg}<16'b0100111111010101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100111111010101)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0100111111010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0100111111010111)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==16'b0100111111011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0100111111011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0100111111011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100111111011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0100111111011100) && ({row_reg, col_reg}<16'b0100111111011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100111111011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100111111100000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0100111111100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0100111111100010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0100111111100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100111111100100) && ({row_reg, col_reg}<16'b0100111111101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100111111101001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0100111111101010) && ({row_reg, col_reg}<16'b0100111111110000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0100111111110000) && ({row_reg, col_reg}<16'b0100111111110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0100111111110111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0100111111111000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100111111111001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0100111111111010) && ({row_reg, col_reg}<16'b0100111111111101)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0100111111111101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0100111111111110)) color_data = 12'b010001010011;

		if(({row_reg, col_reg}==16'b0100111111111111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101000000000000) && ({row_reg, col_reg}<16'b0101000000000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000000000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101000000000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000000000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000000000110) && ({row_reg, col_reg}<16'b0101000000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101000000001010) && ({row_reg, col_reg}<16'b0101000000001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101000000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000000001101) && ({row_reg, col_reg}<16'b0101000000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000000001111) && ({row_reg, col_reg}<16'b0101000000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000000010010) && ({row_reg, col_reg}<16'b0101000000111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101000000111010) && ({row_reg, col_reg}<16'b0101000000111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000000111101) && ({row_reg, col_reg}<16'b0101000001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101000001100011) && ({row_reg, col_reg}<16'b0101000001100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000001100101) && ({row_reg, col_reg}<16'b0101000001100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101000001100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000001101000) && ({row_reg, col_reg}<16'b0101000001101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000001101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000001101011) && ({row_reg, col_reg}<16'b0101000001101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101000001101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000001101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101000001101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000001110000) && ({row_reg, col_reg}<16'b0101000001110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101000001110010) && ({row_reg, col_reg}<16'b0101000001110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000001110101) && ({row_reg, col_reg}<16'b0101000001110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101000001110111) && ({row_reg, col_reg}<16'b0101000001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000001111100) && ({row_reg, col_reg}<16'b0101000001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101000001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000010000001) && ({row_reg, col_reg}<16'b0101000010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101000010010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000010010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000010010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000010010111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000010011000) && ({row_reg, col_reg}<16'b0101000010011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101000010011101) && ({row_reg, col_reg}<16'b0101000010011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000010011111) && ({row_reg, col_reg}<16'b0101000010100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000010100001) && ({row_reg, col_reg}<16'b0101000010100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000010100011) && ({row_reg, col_reg}<16'b0101000010100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101000010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101000010100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000010101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101000010101001) && ({row_reg, col_reg}<16'b0101000010101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000010101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101000010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000010101110) && ({row_reg, col_reg}<16'b0101000010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000010110000) && ({row_reg, col_reg}<16'b0101000010110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101000010110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101000010110011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0101000010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000010110101) && ({row_reg, col_reg}<16'b0101000010110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101000010110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101000010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000010111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000010111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101000010111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101000010111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000010111110) && ({row_reg, col_reg}<16'b0101000011000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000011000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000011000010) && ({row_reg, col_reg}<16'b0101000011000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101000011000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000011000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000011001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000011001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101000011001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000011001011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101000011001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101000011001101) && ({row_reg, col_reg}<16'b0101000011010010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101000011010010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101000011010011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101000011010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101000011010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000011010110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101000011010111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101000011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101000011011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101000011011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101000011011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000011011100) && ({row_reg, col_reg}<16'b0101000011011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101000011011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101000011100000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101000011100001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000011100010) && ({row_reg, col_reg}<16'b0101000011100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101000011100100) && ({row_reg, col_reg}<16'b0101000011101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000011101010) && ({row_reg, col_reg}<16'b0101000011110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000011110000) && ({row_reg, col_reg}<16'b0101000011110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000011110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000011110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101000011110101) && ({row_reg, col_reg}<16'b0101000011110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000011110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101000011111000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101000011111001) && ({row_reg, col_reg}<16'b0101000011111011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101000011111011) && ({row_reg, col_reg}<16'b0101000011111110)) color_data = 12'b010001010011;

		if(({row_reg, col_reg}>=16'b0101000011111110) && ({row_reg, col_reg}<16'b0101000100000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101000100000000) && ({row_reg, col_reg}<16'b0101000100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000100000101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101000100000110) && ({row_reg, col_reg}<16'b0101000100001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101000100001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101000100001011) && ({row_reg, col_reg}<16'b0101000100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000100001101) && ({row_reg, col_reg}<16'b0101000100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000100010010) && ({row_reg, col_reg}<16'b0101000100111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101000100111010) && ({row_reg, col_reg}<16'b0101000100111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000100111101) && ({row_reg, col_reg}<16'b0101000100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101000100111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000101000000) && ({row_reg, col_reg}<16'b0101000101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101000101100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101000101100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000101100101) && ({row_reg, col_reg}<16'b0101000101100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101000101100111) && ({row_reg, col_reg}<16'b0101000101101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000101101001) && ({row_reg, col_reg}<16'b0101000101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000101101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000101101101) && ({row_reg, col_reg}<16'b0101000101101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000101101111) && ({row_reg, col_reg}<16'b0101000101110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101000101110111) && ({row_reg, col_reg}<16'b0101000101111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000101111100) && ({row_reg, col_reg}<16'b0101000101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101000101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000110000001) && ({row_reg, col_reg}<16'b0101000110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101000110010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000110010101) && ({row_reg, col_reg}<16'b0101000110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000110010111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000110011000) && ({row_reg, col_reg}<16'b0101000110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101000110011101) && ({row_reg, col_reg}<16'b0101000110011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000110100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101000110100001) && ({row_reg, col_reg}<16'b0101000110100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000110100011) && ({row_reg, col_reg}<16'b0101000110100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101000110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101000110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000110101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101000110101001) && ({row_reg, col_reg}<16'b0101000110101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101000110101110) && ({row_reg, col_reg}<16'b0101000110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000110110000) && ({row_reg, col_reg}<16'b0101000110110100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101000110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000110110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101000110110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000110110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101000110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000110111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000110111011) && ({row_reg, col_reg}<16'b0101000110111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101000110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000110111110) && ({row_reg, col_reg}<16'b0101000111000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101000111000001) && ({row_reg, col_reg}<16'b0101000111000011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000111000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101000111000100) && ({row_reg, col_reg}<16'b0101000111000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000111000110) && ({row_reg, col_reg}<16'b0101000111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000111001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101000111001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000111001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101000111001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101000111001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101000111001110) && ({row_reg, col_reg}<16'b0101000111010000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101000111010000)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0101000111010001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101000111010010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101000111010011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101000111010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101000111010101) && ({row_reg, col_reg}<16'b0101000111010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000111010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000111011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101000111011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101000111011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101000111011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000111011100) && ({row_reg, col_reg}<16'b0101000111011111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101000111011111) && ({row_reg, col_reg}<16'b0101000111100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101000111100010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101000111100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101000111100100) && ({row_reg, col_reg}<16'b0101000111101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101000111101100) && ({row_reg, col_reg}<16'b0101000111101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101000111101110) && ({row_reg, col_reg}<16'b0101000111110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000111110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101000111110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101000111110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101000111110101) && ({row_reg, col_reg}<16'b0101000111110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101000111110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101000111111000)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0101000111111001)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0101000111111010) && ({row_reg, col_reg}<16'b0101000111111110)) color_data = 12'b010001010011;

		if(({row_reg, col_reg}>=16'b0101000111111110) && ({row_reg, col_reg}<16'b0101001000000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101001000000000) && ({row_reg, col_reg}<16'b0101001000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001000000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101001000000110) && ({row_reg, col_reg}<16'b0101001000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101001000001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101001000001011) && ({row_reg, col_reg}<16'b0101001000001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001000001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001000001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101001000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001000010010) && ({row_reg, col_reg}<16'b0101001000111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101001000111010) && ({row_reg, col_reg}<16'b0101001000111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001000111101) && ({row_reg, col_reg}<16'b0101001001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101001001100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001001100100) && ({row_reg, col_reg}<16'b0101001001101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001001101010) && ({row_reg, col_reg}<16'b0101001001101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001001101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001001101101) && ({row_reg, col_reg}<16'b0101001001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001001110000) && ({row_reg, col_reg}<16'b0101001001110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101001001110010) && ({row_reg, col_reg}<16'b0101001001110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001001110100) && ({row_reg, col_reg}<16'b0101001001110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101001001110111) && ({row_reg, col_reg}<16'b0101001001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001001111100) && ({row_reg, col_reg}<16'b0101001001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101001001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001010000001) && ({row_reg, col_reg}<16'b0101001010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101001010010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001010010101) && ({row_reg, col_reg}<16'b0101001010010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001010010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001010011000) && ({row_reg, col_reg}<16'b0101001010011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101001010011101) && ({row_reg, col_reg}<16'b0101001010011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101001010011111) && ({row_reg, col_reg}<16'b0101001010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001010100011) && ({row_reg, col_reg}<16'b0101001010100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101001010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001010100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001010101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101001010101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001010101010) && ({row_reg, col_reg}<16'b0101001010110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101001010110011) && ({row_reg, col_reg}<16'b0101001010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101001010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001010110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101001010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001010111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101001010111010) && ({row_reg, col_reg}<16'b0101001010111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001010111100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0101001010111101) && ({row_reg, col_reg}<16'b0101001011000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001011000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101001011000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001011000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101001011000100) && ({row_reg, col_reg}<16'b0101001011000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001011000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001011000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101001011001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001011001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101001011001010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0101001011001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101001011001100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001011001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101001011001110)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}>=16'b0101001011001111) && ({row_reg, col_reg}<16'b0101001011010001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0101001011010001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101001011010010)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==16'b0101001011010011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101001011010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001011010101)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0101001011010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101001011010111) && ({row_reg, col_reg}<16'b0101001011011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101001011011010) && ({row_reg, col_reg}<16'b0101001011011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101001011011100) && ({row_reg, col_reg}<16'b0101001011100000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101001011100000) && ({row_reg, col_reg}<16'b0101001011100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101001011100010) && ({row_reg, col_reg}<16'b0101001011100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001011100110)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}>=16'b0101001011100111) && ({row_reg, col_reg}<16'b0101001011101010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001011101010)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}>=16'b0101001011101011) && ({row_reg, col_reg}<16'b0101001011110001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001011110001)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}>=16'b0101001011110010) && ({row_reg, col_reg}<16'b0101001011110110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001011110110)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}>=16'b0101001011110111) && ({row_reg, col_reg}<16'b0101001011111001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001011111001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101001011111010)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0101001011111011) && ({row_reg, col_reg}<16'b0101001011111101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101001011111101)) color_data = 12'b010001010011;

		if(({row_reg, col_reg}>=16'b0101001011111110) && ({row_reg, col_reg}<16'b0101001100000000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101001100000000) && ({row_reg, col_reg}<16'b0101001100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001100000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101001100000110) && ({row_reg, col_reg}<16'b0101001100001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101001100001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101001100001011) && ({row_reg, col_reg}<16'b0101001100001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001100001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001100001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101001100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001100010010) && ({row_reg, col_reg}<16'b0101001100111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101001100111010) && ({row_reg, col_reg}<16'b0101001100111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001100111101) && ({row_reg, col_reg}<16'b0101001101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101001101100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001101100100) && ({row_reg, col_reg}<16'b0101001101101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001101101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001101101101) && ({row_reg, col_reg}<16'b0101001101110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001101110101) && ({row_reg, col_reg}<16'b0101001101110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101001101110111) && ({row_reg, col_reg}<16'b0101001101111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001101111101) && ({row_reg, col_reg}<16'b0101001101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101001101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101001110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101001110000001) && ({row_reg, col_reg}<16'b0101001110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101001110010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001110010101) && ({row_reg, col_reg}<16'b0101001110011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101001110011000) && ({row_reg, col_reg}<16'b0101001110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101001110011101) && ({row_reg, col_reg}<16'b0101001110100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001110100000) && ({row_reg, col_reg}<16'b0101001110100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101001110100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001110100011) && ({row_reg, col_reg}<16'b0101001110100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101001110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101001110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001110101010) && ({row_reg, col_reg}<16'b0101001110110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001110110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101001110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101001110110110) && ({row_reg, col_reg}<16'b0101001110111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101001110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101001110111001) && ({row_reg, col_reg}<16'b0101001110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101001110111011) && ({row_reg, col_reg}<16'b0101001110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101001110111110) && ({row_reg, col_reg}<16'b0101001111000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101001111000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001111000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101001111000100) && ({row_reg, col_reg}<16'b0101001111000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101001111000110) && ({row_reg, col_reg}<16'b0101001111001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101001111001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101001111001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101001111001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101001111001100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101001111001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101001111001110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101001111001111)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}>=16'b0101001111010000) && ({row_reg, col_reg}<16'b0101001111010010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101001111010010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101001111010011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101001111010100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101001111010101) && ({row_reg, col_reg}<16'b0101001111010111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101001111010111) && ({row_reg, col_reg}<16'b0101001111011010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0101001111011010) && ({row_reg, col_reg}<16'b0101001111100110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101001111100110) && ({row_reg, col_reg}<16'b0101001111101101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101001111101101) && ({row_reg, col_reg}<16'b0101001111110000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101001111110000) && ({row_reg, col_reg}<16'b0101001111110010)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0101001111110010) && ({row_reg, col_reg}<16'b0101001111110101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101001111110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101001111110110)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101001111110111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101001111111000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101001111111001)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==16'b0101001111111010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101001111111011)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}>=16'b0101001111111100) && ({row_reg, col_reg}<16'b0101001111111110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101001111111110)) color_data = 12'b010101000011;

		if(({row_reg, col_reg}==16'b0101001111111111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101010000000000) && ({row_reg, col_reg}<16'b0101010000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010000000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101010000000110) && ({row_reg, col_reg}<16'b0101010000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101010000001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101010000001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010000001101) && ({row_reg, col_reg}<16'b0101010000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010000001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101010000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010000010010) && ({row_reg, col_reg}<16'b0101010000110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101010000110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010000110100) && ({row_reg, col_reg}<16'b0101010000111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101010000111010) && ({row_reg, col_reg}<16'b0101010000111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010000111101) && ({row_reg, col_reg}<16'b0101010001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101010001100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010001100100) && ({row_reg, col_reg}<16'b0101010001101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010001101011) && ({row_reg, col_reg}<16'b0101010001101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010001101101) && ({row_reg, col_reg}<16'b0101010001110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010001110000) && ({row_reg, col_reg}<16'b0101010001110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010001110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010001110100) && ({row_reg, col_reg}<16'b0101010001110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010001110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101010001110111) && ({row_reg, col_reg}<16'b0101010010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010010000001) && ({row_reg, col_reg}<16'b0101010010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101010010010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010010010101) && ({row_reg, col_reg}<16'b0101010010011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010010011000) && ({row_reg, col_reg}<16'b0101010010011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101010010011101) && ({row_reg, col_reg}<16'b0101010010011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010010011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101010010100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101010010100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101010010100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010010100011) && ({row_reg, col_reg}<16'b0101010010100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101010010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101010010100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101010010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101010010101001) && ({row_reg, col_reg}<16'b0101010010101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010010101011) && ({row_reg, col_reg}<16'b0101010010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010010110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101010010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010010110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101010010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101010010110110) && ({row_reg, col_reg}<16'b0101010010111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101010010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101010010111001) && ({row_reg, col_reg}<16'b0101010010111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101010010111011) && ({row_reg, col_reg}<16'b0101010010111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101010010111101) && ({row_reg, col_reg}<16'b0101010011000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101010011000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101010011000010) && ({row_reg, col_reg}<16'b0101010011000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101010011000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010011000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010011000110) && ({row_reg, col_reg}<16'b0101010011001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101010011001001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==16'b0101010011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010011001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101010011001100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0101010011001101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101010011001110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010011001111)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0101010011010000) && ({row_reg, col_reg}<16'b0101010011010010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101010011010010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101010011010011) && ({row_reg, col_reg}<16'b0101010011010111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010011010111)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101010011011000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101010011011001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101010011011010) && ({row_reg, col_reg}<16'b0101010011100011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010011100011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101010011100100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101010011100101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101010011100110) && ({row_reg, col_reg}<16'b0101010011101101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010011101101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101010011101110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101010011101111)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0101010011110000) && ({row_reg, col_reg}<16'b0101010011110010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010011110010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101010011110011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101010011110100)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0101010011110101) && ({row_reg, col_reg}<16'b0101010011111000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010011111000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101010011111001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101010011111010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101010011111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101010011111100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101010011111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101010011111110)) color_data = 12'b010101000011;

		if(({row_reg, col_reg}==16'b0101010011111111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101010100000000) && ({row_reg, col_reg}<16'b0101010100000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010100000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010100000011) && ({row_reg, col_reg}<16'b0101010100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010100000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101010100000110) && ({row_reg, col_reg}<16'b0101010100001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101010100001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101010100001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010100001101) && ({row_reg, col_reg}<16'b0101010100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010100010010) && ({row_reg, col_reg}<16'b0101010100111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101010100111010) && ({row_reg, col_reg}<16'b0101010100111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010100111101) && ({row_reg, col_reg}<16'b0101010101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101010101100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010101100100) && ({row_reg, col_reg}<16'b0101010101101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010101101011) && ({row_reg, col_reg}<16'b0101010101101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010101101101) && ({row_reg, col_reg}<16'b0101010101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010101101111) && ({row_reg, col_reg}<16'b0101010110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010110000010) && ({row_reg, col_reg}<16'b0101010110010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101010110010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101010110010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010110010101) && ({row_reg, col_reg}<16'b0101010110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010110010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010110011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010110011001) && ({row_reg, col_reg}<16'b0101010110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101010110011101) && ({row_reg, col_reg}<16'b0101010110011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010110100000) && ({row_reg, col_reg}<16'b0101010110100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101010110100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101010110100011) && ({row_reg, col_reg}<16'b0101010110100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101010110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010110100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101010110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101010110101001) && ({row_reg, col_reg}<16'b0101010110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010110101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101010110101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101010110101101) && ({row_reg, col_reg}<16'b0101010110110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101010110110001) && ({row_reg, col_reg}<16'b0101010110110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101010110110011) && ({row_reg, col_reg}<16'b0101010110110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101010110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101010110110110) && ({row_reg, col_reg}<16'b0101010110111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101010110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101010110111001) && ({row_reg, col_reg}<16'b0101010110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101010110111011) && ({row_reg, col_reg}<16'b0101010110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101010110111101) && ({row_reg, col_reg}<16'b0101010111000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101010111000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101010111000010) && ({row_reg, col_reg}<16'b0101010111000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101010111000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101010111000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101010111000110) && ({row_reg, col_reg}<16'b0101010111001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101010111001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101010111001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101010111001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010111001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101010111001101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101010111001110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010111001111)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101010111010000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101010111010001)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0101010111010010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101010111010011) && ({row_reg, col_reg}<16'b0101010111010101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101010111010101) && ({row_reg, col_reg}<16'b0101010111010111)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0101010111010111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101010111011000)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0101010111011001)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0101010111011010) && ({row_reg, col_reg}<16'b0101010111011101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010111011101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101010111011110) && ({row_reg, col_reg}<16'b0101010111100011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010111100011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101010111100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101010111100101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010111100110)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}>=16'b0101010111100111) && ({row_reg, col_reg}<16'b0101010111101011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010111101011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101010111101100) && ({row_reg, col_reg}<16'b0101010111101110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101010111101110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101010111101111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101010111110000) && ({row_reg, col_reg}<16'b0101010111110011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101010111110011) && ({row_reg, col_reg}<16'b0101010111110111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101010111110111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101010111111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101010111111001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101010111111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101010111111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101010111111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101010111111101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101010111111110)) color_data = 12'b010101000011;

		if(({row_reg, col_reg}==16'b0101010111111111)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0101011000000000) && ({row_reg, col_reg}<16'b0101011000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011000000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101011000000110) && ({row_reg, col_reg}<16'b0101011000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101011000001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101011000001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011000001101) && ({row_reg, col_reg}<16'b0101011000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011000010010) && ({row_reg, col_reg}<16'b0101011000111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011000111010) && ({row_reg, col_reg}<16'b0101011000111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011000111101) && ({row_reg, col_reg}<16'b0101011001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101011001100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011001100100) && ({row_reg, col_reg}<16'b0101011001101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011001101011) && ({row_reg, col_reg}<16'b0101011001101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011001101101) && ({row_reg, col_reg}<16'b0101011001101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011001101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101011001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011001110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011001110010) && ({row_reg, col_reg}<16'b0101011010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011010000010) && ({row_reg, col_reg}<16'b0101011010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011010010100) && ({row_reg, col_reg}<16'b0101011010010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011010010110) && ({row_reg, col_reg}<16'b0101011010011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011010011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011010011001) && ({row_reg, col_reg}<16'b0101011010011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011010011101) && ({row_reg, col_reg}<16'b0101011010100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011010100000) && ({row_reg, col_reg}<16'b0101011010100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101011010100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011010100011) && ({row_reg, col_reg}<16'b0101011010100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101011010100101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0101011010100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101011010100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011010101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101011010101001) && ({row_reg, col_reg}<16'b0101011010101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011010101011) && ({row_reg, col_reg}<16'b0101011010101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101011010101101) && ({row_reg, col_reg}<16'b0101011010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101011010110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101011010110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101011010110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101011010110011) && ({row_reg, col_reg}<16'b0101011010110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101011010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101011010110110) && ({row_reg, col_reg}<16'b0101011010111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101011010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101011010111001) && ({row_reg, col_reg}<16'b0101011010111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101011010111011) && ({row_reg, col_reg}<16'b0101011010111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101011010111101) && ({row_reg, col_reg}<16'b0101011011000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101011011000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011011000010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101011011000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101011011000100) && ({row_reg, col_reg}<16'b0101011011000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011011000110) && ({row_reg, col_reg}<16'b0101011011001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101011011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101011011001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011011001100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101011011001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101011011001110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011011001111)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0101011011010000) && ({row_reg, col_reg}<16'b0101011011010010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101011011010010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101011011010011) && ({row_reg, col_reg}<16'b0101011011010111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011011010111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101011011011000) && ({row_reg, col_reg}<16'b0101011011011010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101011011011010)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0101011011011011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011011011100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101011011011101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101011011011110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101011011011111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101011011100000) && ({row_reg, col_reg}<16'b0101011011100010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101011011100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011011100011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101011011100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101011011100101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101011011100110) && ({row_reg, col_reg}<16'b0101011011101010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011011101010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101011011101011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101011011101100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101011011101101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0101011011101110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011011101111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101011011110000) && ({row_reg, col_reg}<16'b0101011011110011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101011011110011) && ({row_reg, col_reg}<16'b0101011011110110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011011110110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101011011110111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101011011111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101011011111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101011011111010) && ({row_reg, col_reg}<16'b0101011011111100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101011011111100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0101011011111101) && ({row_reg, col_reg}<16'b0101011011111111)) color_data = 12'b010101000011;

		if(({row_reg, col_reg}==16'b0101011011111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101011100000000) && ({row_reg, col_reg}<16'b0101011100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011100000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101011100000110) && ({row_reg, col_reg}<16'b0101011100001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101011100001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101011100001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011100001101) && ({row_reg, col_reg}<16'b0101011100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011100010010) && ({row_reg, col_reg}<16'b0101011100111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011100111011) && ({row_reg, col_reg}<16'b0101011100111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011100111101) && ({row_reg, col_reg}<16'b0101011101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101011101100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011101100100) && ({row_reg, col_reg}<16'b0101011101101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011101101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101011101101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011101101010) && ({row_reg, col_reg}<16'b0101011101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011101101100) && ({row_reg, col_reg}<16'b0101011101101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011101101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101011101110000) && ({row_reg, col_reg}<16'b0101011101111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011101111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011101111110) && ({row_reg, col_reg}<16'b0101011110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011110000001) && ({row_reg, col_reg}<16'b0101011110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101011110010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011110010101) && ({row_reg, col_reg}<16'b0101011110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011110010111) && ({row_reg, col_reg}<16'b0101011110011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101011110011001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011110011010) && ({row_reg, col_reg}<16'b0101011110011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011110011100) && ({row_reg, col_reg}<16'b0101011110100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011110100000) && ({row_reg, col_reg}<16'b0101011110100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101011110100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011110100011) && ({row_reg, col_reg}<16'b0101011110100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101011110100110) && ({row_reg, col_reg}<16'b0101011110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101011110101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101011110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011110101011) && ({row_reg, col_reg}<16'b0101011110101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101011110101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101011110101110) && ({row_reg, col_reg}<16'b0101011110110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101011110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101011110110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101011110110101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0101011110110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101011110110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101011110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101011110111001) && ({row_reg, col_reg}<16'b0101011110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101011110111011) && ({row_reg, col_reg}<16'b0101011110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101011110111110) && ({row_reg, col_reg}<16'b0101011111000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101011111000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101011111000011) && ({row_reg, col_reg}<16'b0101011111000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101011111000101) && ({row_reg, col_reg}<16'b0101011111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101011111000111) && ({row_reg, col_reg}<16'b0101011111001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101011111001001) && ({row_reg, col_reg}<16'b0101011111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101011111001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101011111001100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0101011111001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101011111001110)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101011111001111) && ({row_reg, col_reg}<16'b0101011111010001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101011111010001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101011111010010) && ({row_reg, col_reg}<16'b0101011111010100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011111010100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0101011111010101) && ({row_reg, col_reg}<16'b0101011111010111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101011111010111)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0101011111011000) && ({row_reg, col_reg}<16'b0101011111011010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011111011010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101011111011011) && ({row_reg, col_reg}<16'b0101011111011101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101011111011101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101011111011110) && ({row_reg, col_reg}<16'b0101011111100000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101011111100000) && ({row_reg, col_reg}<16'b0101011111100010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101011111100010) && ({row_reg, col_reg}<16'b0101011111100100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011111100100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101011111100101) && ({row_reg, col_reg}<16'b0101011111100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101011111100111) && ({row_reg, col_reg}<16'b0101011111101001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011111101001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101011111101010)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101011111101011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101011111101100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101011111101101) && ({row_reg, col_reg}<16'b0101011111101111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101011111101111)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0101011111110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101011111110001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0101011111110010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101011111110011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101011111110100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101011111110101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101011111110110) && ({row_reg, col_reg}<16'b0101011111111000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101011111111000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101011111111001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101011111111010)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101011111111011) && ({row_reg, col_reg}<16'b0101011111111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101011111111101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101011111111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0101011111111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101100000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100000000001) && ({row_reg, col_reg}<16'b0101100000000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100000000011) && ({row_reg, col_reg}<16'b0101100000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100000000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101100000000110) && ({row_reg, col_reg}<16'b0101100000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101100000001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101100000001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100000001101) && ({row_reg, col_reg}<16'b0101100000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100000010001) && ({row_reg, col_reg}<16'b0101100001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100001100011) && ({row_reg, col_reg}<16'b0101100001101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100001101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100001101011) && ({row_reg, col_reg}<16'b0101100001101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100001101101) && ({row_reg, col_reg}<16'b0101100001101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100001101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101100001110000) && ({row_reg, col_reg}<16'b0101100001110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100001110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101100001110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100001110110) && ({row_reg, col_reg}<16'b0101100001111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100001111000) && ({row_reg, col_reg}<16'b0101100001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100001111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101100001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100001111110) && ({row_reg, col_reg}<16'b0101100010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100010000001) && ({row_reg, col_reg}<16'b0101100010010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100010010101) && ({row_reg, col_reg}<16'b0101100010011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100010011000) && ({row_reg, col_reg}<16'b0101100010100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100010100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101100010100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100010100010) && ({row_reg, col_reg}<16'b0101100010100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100010100101) && ({row_reg, col_reg}<16'b0101100010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101100010101001) && ({row_reg, col_reg}<16'b0101100010101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100010101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101100010101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101100010101101) && ({row_reg, col_reg}<16'b0101100010101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100010101111) && ({row_reg, col_reg}<16'b0101100010110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101100010110011) && ({row_reg, col_reg}<16'b0101100010110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101100010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100010110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101100010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101100010111001) && ({row_reg, col_reg}<16'b0101100010111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101100010111011) && ({row_reg, col_reg}<16'b0101100010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101100010111110) && ({row_reg, col_reg}<16'b0101100011000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101100011000010) && ({row_reg, col_reg}<16'b0101100011000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101100011000100) && ({row_reg, col_reg}<16'b0101100011000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101100011000110) && ({row_reg, col_reg}<16'b0101100011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100011001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100011001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101100011001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101100011001100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101100011001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101100011001110)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==16'b0101100011001111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101100011010000)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101100011010001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0101100011010010) && ({row_reg, col_reg}<16'b0101100011010100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101100011010100) && ({row_reg, col_reg}<16'b0101100011010111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101100011010111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101100011011000) && ({row_reg, col_reg}<16'b0101100011011011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101100011011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101100011011100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0101100011011101) && ({row_reg, col_reg}<16'b0101100011100000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101100011100000) && ({row_reg, col_reg}<16'b0101100011100010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101100011100010) && ({row_reg, col_reg}<16'b0101100011100101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101100011100101) && ({row_reg, col_reg}<16'b0101100011100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101100011100111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101100011101000)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101100011101001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101100011101010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101100011101011) && ({row_reg, col_reg}<16'b0101100011101111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101100011101111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101100011110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101100011110001) && ({row_reg, col_reg}<16'b0101100011110011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101100011110011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101100011110100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101100011110101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101100011110110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101100011110111)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=16'b0101100011111000) && ({row_reg, col_reg}<16'b0101100011111010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101100011111010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101100011111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101100011111100) && ({row_reg, col_reg}<16'b0101100011111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101100011111110)) color_data = 12'b001100110010;

		if(({row_reg, col_reg}==16'b0101100011111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100100000001) && ({row_reg, col_reg}<16'b0101100100000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100100000011) && ({row_reg, col_reg}<16'b0101100100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100100000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101100100000110) && ({row_reg, col_reg}<16'b0101100100001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101100100001010) && ({row_reg, col_reg}<16'b0101100100001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101100100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100100001101) && ({row_reg, col_reg}<16'b0101100100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100100001111) && ({row_reg, col_reg}<16'b0101100100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100100010001) && ({row_reg, col_reg}<16'b0101100100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101100100110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100100110100) && ({row_reg, col_reg}<16'b0101100101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101100101100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100101100011) && ({row_reg, col_reg}<16'b0101100101101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100101101000) && ({row_reg, col_reg}<16'b0101100101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100101101011) && ({row_reg, col_reg}<16'b0101100101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101100101101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101100101101110) && ({row_reg, col_reg}<16'b0101100101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100101110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101100101110001) && ({row_reg, col_reg}<16'b0101100101110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100101110110) && ({row_reg, col_reg}<16'b0101100101111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100101111001) && ({row_reg, col_reg}<16'b0101100101111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100101111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101100101111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100101111110) && ({row_reg, col_reg}<16'b0101100110000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101100110000001) && ({row_reg, col_reg}<16'b0101100110010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100110010101) && ({row_reg, col_reg}<16'b0101100110011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100110011000) && ({row_reg, col_reg}<16'b0101100110011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100110011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100110011011) && ({row_reg, col_reg}<16'b0101100110100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100110100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101100110100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100110100010) && ({row_reg, col_reg}<16'b0101100110100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100110100110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0101100110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101100110101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100110101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101100110101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100110101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101100110101101) && ({row_reg, col_reg}<16'b0101100110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101100110110000) && ({row_reg, col_reg}<16'b0101100110110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101100110110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101100110110011) && ({row_reg, col_reg}<16'b0101100110110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101100110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101100110110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100110110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101100110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101100110111001) && ({row_reg, col_reg}<16'b0101100110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101100110111011) && ({row_reg, col_reg}<16'b0101100110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101100110111110) && ({row_reg, col_reg}<16'b0101100111000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101100111000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100111000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101100111000110) && ({row_reg, col_reg}<16'b0101100111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101100111001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101100111001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101100111001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101100111001100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101100111001101)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}>=16'b0101100111001110) && ({row_reg, col_reg}<16'b0101100111010000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101100111010000) && ({row_reg, col_reg}<16'b0101100111010010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101100111010010)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101100111010011)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0101100111010100) && ({row_reg, col_reg}<16'b0101100111100000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101100111100000) && ({row_reg, col_reg}<16'b0101100111100010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101100111100010) && ({row_reg, col_reg}<16'b0101100111101001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101100111101001)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101100111101010) && ({row_reg, col_reg}<16'b0101100111111011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101100111111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101100111111100) && ({row_reg, col_reg}<16'b0101100111111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101100111111110)) color_data = 12'b001100110010;

		if(({row_reg, col_reg}==16'b0101100111111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101101000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101000000001) && ({row_reg, col_reg}<16'b0101101000000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101000000011) && ({row_reg, col_reg}<16'b0101101000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101000000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101101000000110) && ({row_reg, col_reg}<16'b0101101000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101101000001001) && ({row_reg, col_reg}<16'b0101101000001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101101000001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101000001101) && ({row_reg, col_reg}<16'b0101101000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101000001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101000010001) && ({row_reg, col_reg}<16'b0101101001100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101101001100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101001100011) && ({row_reg, col_reg}<16'b0101101001101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101001101000) && ({row_reg, col_reg}<16'b0101101001101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101001101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101001101011) && ({row_reg, col_reg}<16'b0101101001101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101101001101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101101001101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101001101111) && ({row_reg, col_reg}<16'b0101101001110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101101001110010) && ({row_reg, col_reg}<16'b0101101001110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101001110110) && ({row_reg, col_reg}<16'b0101101001111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101001111000) && ({row_reg, col_reg}<16'b0101101001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101001111100) && ({row_reg, col_reg}<16'b0101101001111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101101001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101001111111) && ({row_reg, col_reg}<16'b0101101010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101010000001) && ({row_reg, col_reg}<16'b0101101010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101101010010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101010010101) && ({row_reg, col_reg}<16'b0101101010011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101010011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101010011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101010011101) && ({row_reg, col_reg}<16'b0101101010100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101010100000) && ({row_reg, col_reg}<16'b0101101010100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101101010100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101010100011) && ({row_reg, col_reg}<16'b0101101010100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101010100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101101010100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101101010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101101010101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101010101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101101010101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101010101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101101010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101010101110) && ({row_reg, col_reg}<16'b0101101010110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101010110001) && ({row_reg, col_reg}<16'b0101101010110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101101010110011) && ({row_reg, col_reg}<16'b0101101010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101101010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101010110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101010111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101101010111011) && ({row_reg, col_reg}<16'b0101101010111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101101010111101) && ({row_reg, col_reg}<16'b0101101011000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101011000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101101011000011) && ({row_reg, col_reg}<16'b0101101011000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101011000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101101011000110) && ({row_reg, col_reg}<16'b0101101011001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101101011001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101011001001) && ({row_reg, col_reg}<16'b0101101011001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101101011001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101011001100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101101011001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101101011001110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101101011001111)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0101101011010000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101101011010001)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0101101011010010) && ({row_reg, col_reg}<16'b0101101011010100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101101011010100)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101101011010101) && ({row_reg, col_reg}<16'b0101101011100000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101101011100000) && ({row_reg, col_reg}<16'b0101101011100010)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}>=16'b0101101011100010) && ({row_reg, col_reg}<16'b0101101011101000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101101011101000)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0101101011101001)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0101101011101010)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0101101011101011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101101011101100) && ({row_reg, col_reg}<16'b0101101011101110)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=16'b0101101011101110) && ({row_reg, col_reg}<16'b0101101011111100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101101011111100) && ({row_reg, col_reg}<16'b0101101011111110)) color_data = 12'b010101000011;

		if(({row_reg, col_reg}>=16'b0101101011111110) && ({row_reg, col_reg}<16'b0101101100000000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=16'b0101101100000000) && ({row_reg, col_reg}<16'b0101101100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101100000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101101100000110) && ({row_reg, col_reg}<16'b0101101100001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101101100001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101101100001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101100001101) && ({row_reg, col_reg}<16'b0101101100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101100001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101101100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101100010010) && ({row_reg, col_reg}<16'b0101101101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101101101100011) && ({row_reg, col_reg}<16'b0101101101101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101101101000) && ({row_reg, col_reg}<16'b0101101101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101101101011) && ({row_reg, col_reg}<16'b0101101101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101101101101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101101101110) && ({row_reg, col_reg}<16'b0101101101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101101110000) && ({row_reg, col_reg}<16'b0101101101110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101101101110010) && ({row_reg, col_reg}<16'b0101101101110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101101110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101101101110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101101110111) && ({row_reg, col_reg}<16'b0101101101111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101101111100) && ({row_reg, col_reg}<16'b0101101101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101101101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101101111111) && ({row_reg, col_reg}<16'b0101101110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101110000010) && ({row_reg, col_reg}<16'b0101101110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101101110010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101110010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101110010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101110010111) && ({row_reg, col_reg}<16'b0101101110011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101101110011011) && ({row_reg, col_reg}<16'b0101101110011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101101110011101) && ({row_reg, col_reg}<16'b0101101110100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101110100000) && ({row_reg, col_reg}<16'b0101101110100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101101110100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101101110100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101101110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101110100110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0101101110100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101101110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101101110101001) && ({row_reg, col_reg}<16'b0101101110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101110101011) && ({row_reg, col_reg}<16'b0101101110101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101101110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101101110101110) && ({row_reg, col_reg}<16'b0101101110110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101110110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101101110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101101110110101) && ({row_reg, col_reg}<16'b0101101110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101101110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101110111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101101110111011) && ({row_reg, col_reg}<16'b0101101110111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101101110111101) && ({row_reg, col_reg}<16'b0101101110111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101101110111111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101101111000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101101111000001) && ({row_reg, col_reg}<16'b0101101111000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101101111000100) && ({row_reg, col_reg}<16'b0101101111000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101101111000110) && ({row_reg, col_reg}<16'b0101101111001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101101111001000) && ({row_reg, col_reg}<16'b0101101111001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101101111001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101101111001011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0101101111001100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0101101111001101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0101101111001110) && ({row_reg, col_reg}<16'b0101101111010000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101101111010000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101101111010001) && ({row_reg, col_reg}<16'b0101101111010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101101111010100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101101111010101)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=16'b0101101111010110) && ({row_reg, col_reg}<16'b0101101111011110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101101111011110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101101111011111)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}>=16'b0101101111100000) && ({row_reg, col_reg}<16'b0101101111100010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0101101111100010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101101111100011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101101111100100) && ({row_reg, col_reg}<16'b0101101111100111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101101111100111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101101111101000)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0101101111101001)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==16'b0101101111101010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0101101111101011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101101111101100) && ({row_reg, col_reg}<16'b0101101111101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==16'b0101101111101110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101101111101111)) color_data = 12'b011001010011;

		if(({row_reg, col_reg}>=16'b0101101111110000) && ({row_reg, col_reg}<16'b0101110000000000)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101110000000000) && ({row_reg, col_reg}<16'b0101110000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110000000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110000000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101110000001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101110000001010) && ({row_reg, col_reg}<16'b0101110000001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110000001101) && ({row_reg, col_reg}<16'b0101110000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110000001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101110000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110000010010) && ({row_reg, col_reg}<16'b0101110001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101110001100011) && ({row_reg, col_reg}<16'b0101110001101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110001101000) && ({row_reg, col_reg}<16'b0101110001101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110001101011) && ({row_reg, col_reg}<16'b0101110001101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101110001101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110001101110) && ({row_reg, col_reg}<16'b0101110001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110001110000) && ({row_reg, col_reg}<16'b0101110001110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101110001110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110001110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110001110111) && ({row_reg, col_reg}<16'b0101110001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110001111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101110001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101110001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110001111111) && ({row_reg, col_reg}<16'b0101110010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110010000010) && ({row_reg, col_reg}<16'b0101110010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101110010010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110010010101) && ({row_reg, col_reg}<16'b0101110010011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101110010011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110010011011) && ({row_reg, col_reg}<16'b0101110010011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110010011101) && ({row_reg, col_reg}<16'b0101110010100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110010100000) && ({row_reg, col_reg}<16'b0101110010100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101110010100011) && ({row_reg, col_reg}<16'b0101110010100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110010100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101110010100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101110010101001) && ({row_reg, col_reg}<16'b0101110010101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101110010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110010101110) && ({row_reg, col_reg}<16'b0101110010110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101110010110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101110010110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110010110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101110010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110010110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101110010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110010111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101110010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110010111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101110010111100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0101110010111101) && ({row_reg, col_reg}<16'b0101110010111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101110010111111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101110011000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101110011000001) && ({row_reg, col_reg}<16'b0101110011000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110011000100) && ({row_reg, col_reg}<16'b0101110011001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101110011001000) && ({row_reg, col_reg}<16'b0101110011001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110011001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101110011001011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0101110011001100)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101110011001101)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101110011001110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101110011001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101110011010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101110011010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101110011010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110011010011) && ({row_reg, col_reg}<16'b0101110011010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101110011010101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101110011010110)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101110011010111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101110011011000)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}>=16'b0101110011011001) && ({row_reg, col_reg}<16'b0101110011011011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101110011011011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101110011011100)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==16'b0101110011011101)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}>=16'b0101110011011110) && ({row_reg, col_reg}<16'b0101110011100000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101110011100000)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0101110011100001)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0101110011100010)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0101110011100011)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}>=16'b0101110011100100) && ({row_reg, col_reg}<16'b0101110011100110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101110011100110) && ({row_reg, col_reg}<16'b0101110011101000)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==16'b0101110011101000)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==16'b0101110011101001)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}>=16'b0101110011101010) && ({row_reg, col_reg}<16'b0101110011101100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101110011101100)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==16'b0101110011101101)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==16'b0101110011101110)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0101110011101111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101110011110000) && ({row_reg, col_reg}<16'b0101110011110100)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==16'b0101110011110100)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101110011110101)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}>=16'b0101110011110110) && ({row_reg, col_reg}<16'b0101110011111001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==16'b0101110011111001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0101110011111010)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101110011111011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101110011111100) && ({row_reg, col_reg}<16'b0101110011111111)) color_data = 12'b011101100100;

		if(({row_reg, col_reg}==16'b0101110011111111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}>=16'b0101110100000000) && ({row_reg, col_reg}<16'b0101110100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110100000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110100000111) && ({row_reg, col_reg}<16'b0101110100001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101110100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101110100001010) && ({row_reg, col_reg}<16'b0101110100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110100001101) && ({row_reg, col_reg}<16'b0101110100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110100001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101110100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110100010010) && ({row_reg, col_reg}<16'b0101110101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101110101100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110101100100) && ({row_reg, col_reg}<16'b0101110101101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110101101000) && ({row_reg, col_reg}<16'b0101110101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110101101011) && ({row_reg, col_reg}<16'b0101110101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101110101101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110101101110) && ({row_reg, col_reg}<16'b0101110101110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110101110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101110101110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110101110100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101110101110101) && ({row_reg, col_reg}<16'b0101110101111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110101111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101110101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110101111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101110101111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101110101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101110101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101110110000001) && ({row_reg, col_reg}<16'b0101110110010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101110110010101) && ({row_reg, col_reg}<16'b0101110110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101110110010111) && ({row_reg, col_reg}<16'b0101110110011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110110011011) && ({row_reg, col_reg}<16'b0101110110011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101110110011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110110011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101110110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110110100000) && ({row_reg, col_reg}<16'b0101110110100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101110110100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101110110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101110110100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101110110100110) && ({row_reg, col_reg}<16'b0101110110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110110101000) && ({row_reg, col_reg}<16'b0101110110101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101110110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101110110101110) && ({row_reg, col_reg}<16'b0101110110110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101110110110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101110110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110110110101) && ({row_reg, col_reg}<16'b0101110110111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101110110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110110111001) && ({row_reg, col_reg}<16'b0101110110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101110110111011) && ({row_reg, col_reg}<16'b0101110110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110110111110) && ({row_reg, col_reg}<16'b0101110111000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101110111000010) && ({row_reg, col_reg}<16'b0101110111000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101110111000110) && ({row_reg, col_reg}<16'b0101110111001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101110111001011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0101110111001100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101110111001101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101110111001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101110111001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101110111010000) && ({row_reg, col_reg}<16'b0101110111010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110111010010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101110111010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101110111010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101110111010101) && ({row_reg, col_reg}<16'b0101110111010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101110111010111) && ({row_reg, col_reg}<16'b0101110111011001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101110111011001) && ({row_reg, col_reg}<16'b0101110111011011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101110111011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101110111011100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101110111011101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101110111011110) && ({row_reg, col_reg}<16'b0101110111100000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101110111100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101110111100001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101110111100010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101110111100011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==16'b0101110111100100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101110111100101) && ({row_reg, col_reg}<16'b0101110111101001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==16'b0101110111101001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101110111101010) && ({row_reg, col_reg}<16'b0101110111101100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0101110111101100) && ({row_reg, col_reg}<16'b0101110111101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101110111101111)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}>=16'b0101110111110000) && ({row_reg, col_reg}<16'b0101110111110010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101110111110010) && ({row_reg, col_reg}<16'b0101110111110100)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101110111110100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101110111110101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0101110111110110) && ({row_reg, col_reg}<16'b0101110111111001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101110111111001) && ({row_reg, col_reg}<16'b0101110111111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0101110111111011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0101110111111100)) color_data = 12'b010101010011;
		if(({row_reg, col_reg}==16'b0101110111111101)) color_data = 12'b011001010011;

		if(({row_reg, col_reg}>=16'b0101110111111110) && ({row_reg, col_reg}<16'b0101111000000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0101111000000000) && ({row_reg, col_reg}<16'b0101111000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111000000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101111000000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111000000111) && ({row_reg, col_reg}<16'b0101111000001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101111000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111000001010) && ({row_reg, col_reg}<16'b0101111000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101111000001100) && ({row_reg, col_reg}<16'b0101111000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111000010010) && ({row_reg, col_reg}<16'b0101111001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111001100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111001100100) && ({row_reg, col_reg}<16'b0101111001101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111001101000) && ({row_reg, col_reg}<16'b0101111001101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101111001101011) && ({row_reg, col_reg}<16'b0101111001101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111001101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111001101110) && ({row_reg, col_reg}<16'b0101111001111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111001111010) && ({row_reg, col_reg}<16'b0101111001111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111001111100) && ({row_reg, col_reg}<16'b0101111001111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101111001111110) && ({row_reg, col_reg}<16'b0101111010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111010000001) && ({row_reg, col_reg}<16'b0101111010010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111010010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111010010110) && ({row_reg, col_reg}<16'b0101111010011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111010011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101111010011001) && ({row_reg, col_reg}<16'b0101111010011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111010011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111010011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111010011101) && ({row_reg, col_reg}<16'b0101111010011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101111010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111010100000) && ({row_reg, col_reg}<16'b0101111010100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111010100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101111010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111010100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101111010100110) && ({row_reg, col_reg}<16'b0101111010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101111010101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101111010101001) && ({row_reg, col_reg}<16'b0101111010101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111010101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101111010101100) && ({row_reg, col_reg}<16'b0101111010101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111010101110) && ({row_reg, col_reg}<16'b0101111010110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0101111010110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101111010110100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0101111010110101) && ({row_reg, col_reg}<16'b0101111010111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101111010111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101111010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111010111011) && ({row_reg, col_reg}<16'b0101111010111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101111010111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111010111110) && ({row_reg, col_reg}<16'b0101111011000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101111011000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101111011000011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0101111011000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0101111011000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111011000110) && ({row_reg, col_reg}<16'b0101111011001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101111011001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111011001001) && ({row_reg, col_reg}<16'b0101111011001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101111011001011) && ({row_reg, col_reg}<16'b0101111011001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101111011001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101111011001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101111011001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101111011010000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0101111011010001) && ({row_reg, col_reg}<16'b0101111011010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111011010101) && ({row_reg, col_reg}<16'b0101111011010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101111011010111) && ({row_reg, col_reg}<16'b0101111011011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0101111011011001) && ({row_reg, col_reg}<16'b0101111011011011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0101111011011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101111011011100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0101111011011101) && ({row_reg, col_reg}<16'b0101111011100000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0101111011100000) && ({row_reg, col_reg}<16'b0101111011100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101111011100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101111011100011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0101111011100100) && ({row_reg, col_reg}<16'b0101111011101001)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0101111011101001) && ({row_reg, col_reg}<16'b0101111011101011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101111011101011)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0101111011101100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0101111011101101) && ({row_reg, col_reg}<16'b0101111011110100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101111011110100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101111011110101)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==16'b0101111011110110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101111011110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101111011111000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101111011111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101111011111010) && ({row_reg, col_reg}<16'b0101111011111100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0101111011111100) && ({row_reg, col_reg}<16'b0101111011111111)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0101111011111111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0101111100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111100000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111100000010) && ({row_reg, col_reg}<16'b0101111100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111100000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101111100000110) && ({row_reg, col_reg}<16'b0101111100001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101111100001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101111100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101111100001100) && ({row_reg, col_reg}<16'b0101111100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111100010010) && ({row_reg, col_reg}<16'b0101111101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111101100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111101100100) && ({row_reg, col_reg}<16'b0101111101101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111101101001) && ({row_reg, col_reg}<16'b0101111101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101111101101011) && ({row_reg, col_reg}<16'b0101111101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111101101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111101101110) && ({row_reg, col_reg}<16'b0101111101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111101111011) && ({row_reg, col_reg}<16'b0101111101111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0101111101111101) && ({row_reg, col_reg}<16'b0101111110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111110000001) && ({row_reg, col_reg}<16'b0101111110010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101111110010101) && ({row_reg, col_reg}<16'b0101111110010111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101111110010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111110011000) && ({row_reg, col_reg}<16'b0101111110011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101111110011010) && ({row_reg, col_reg}<16'b0101111110011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101111110011100) && ({row_reg, col_reg}<16'b0101111110100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111110100000) && ({row_reg, col_reg}<16'b0101111110100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0101111110100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0101111110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111110100101) && ({row_reg, col_reg}<16'b0101111110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111110101000) && ({row_reg, col_reg}<16'b0101111110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111110101011) && ({row_reg, col_reg}<16'b0101111110101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101111110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0101111110101110) && ({row_reg, col_reg}<16'b0101111110110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0101111110110011) && ({row_reg, col_reg}<16'b0101111110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101111110110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0101111110110110) && ({row_reg, col_reg}<16'b0101111110111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0101111110111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0101111110111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111110111010) && ({row_reg, col_reg}<16'b0101111110111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0101111110111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0101111110111101) && ({row_reg, col_reg}<16'b0101111111000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101111111000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0101111111000011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101111111000100)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0101111111000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0101111111000110) && ({row_reg, col_reg}<16'b0101111111001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0101111111001010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0101111111001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0101111111001100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0101111111001101)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0101111111001110) && ({row_reg, col_reg}<16'b0101111111010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0101111111010001) && ({row_reg, col_reg}<16'b0101111111010011)) color_data = 12'b001100100010;

		if(({row_reg, col_reg}>=16'b0101111111010011) && ({row_reg, col_reg}<16'b0110000000000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000000000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000000000010) && ({row_reg, col_reg}<16'b0110000000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000000000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110000000000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110000000000111) && ({row_reg, col_reg}<16'b0110000000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110000000001001) && ({row_reg, col_reg}<16'b0110000000001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110000000001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000000001101) && ({row_reg, col_reg}<16'b0110000000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000000010010) && ({row_reg, col_reg}<16'b0110000001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110000001100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000001100100) && ({row_reg, col_reg}<16'b0110000001101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000001101001) && ({row_reg, col_reg}<16'b0110000001101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000001101011) && ({row_reg, col_reg}<16'b0110000001101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110000001101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000001101110) && ({row_reg, col_reg}<16'b0110000001110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000001110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000001110111) && ({row_reg, col_reg}<16'b0110000001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000001111100) && ({row_reg, col_reg}<16'b0110000001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000001111110) && ({row_reg, col_reg}<16'b0110000010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000010000001) && ({row_reg, col_reg}<16'b0110000010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110000010010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000010010101) && ({row_reg, col_reg}<16'b0110000010011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000010011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000010011010) && ({row_reg, col_reg}<16'b0110000010011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000010011100) && ({row_reg, col_reg}<16'b0110000010100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000010100000) && ({row_reg, col_reg}<16'b0110000010100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110000010100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110000010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000010100101) && ({row_reg, col_reg}<16'b0110000010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110000010101000) && ({row_reg, col_reg}<16'b0110000010101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000010101011) && ({row_reg, col_reg}<16'b0110000010101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110000010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000010101110) && ({row_reg, col_reg}<16'b0110000010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110000010110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110000010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110000010110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000010110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110000010110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000010110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110000010111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110000010111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110000010111010) && ({row_reg, col_reg}<16'b0110000010111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110000010111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110000010111101) && ({row_reg, col_reg}<16'b0110000010111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000010111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110000011000000) && ({row_reg, col_reg}<16'b0110000011000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000011000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110000011000011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0110000011000100)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0110000011000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110000011000110) && ({row_reg, col_reg}<16'b0110000011001011)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}>=16'b0110000011001011) && ({row_reg, col_reg}<16'b0110000100000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110000100000000) && ({row_reg, col_reg}<16'b0110000100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000100000101) && ({row_reg, col_reg}<16'b0110000100000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110000100000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110000100001000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0110000100001001) && ({row_reg, col_reg}<16'b0110000100001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110000100001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000100001101) && ({row_reg, col_reg}<16'b0110000100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000100010001) && ({row_reg, col_reg}<16'b0110000101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110000101100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000101100100) && ({row_reg, col_reg}<16'b0110000101101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000101101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110000101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000101101011) && ({row_reg, col_reg}<16'b0110000101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110000101101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000101101110) && ({row_reg, col_reg}<16'b0110000101110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110000101110111) && ({row_reg, col_reg}<16'b0110000101111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000101111001) && ({row_reg, col_reg}<16'b0110000101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110000101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000101111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110000101111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110000101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000101111111) && ({row_reg, col_reg}<16'b0110000110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000110000010) && ({row_reg, col_reg}<16'b0110000110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110000110010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110000110010101) && ({row_reg, col_reg}<16'b0110000110100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000110100000) && ({row_reg, col_reg}<16'b0110000110100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110000110100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110000110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000110100101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0110000110100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110000110101000) && ({row_reg, col_reg}<16'b0110000110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000110101011) && ({row_reg, col_reg}<16'b0110000110101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110000110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110000110101110) && ({row_reg, col_reg}<16'b0110000110110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110000110110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110000110110011) && ({row_reg, col_reg}<16'b0110000110110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110000110110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110000110110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110000110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110000110111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110000110111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110000110111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110000110111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110000110111110) && ({row_reg, col_reg}<16'b0110000111000000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110000111000000) && ({row_reg, col_reg}<16'b0110000111000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110000111000100) && ({row_reg, col_reg}<16'b0110000111000110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110000111000110) && ({row_reg, col_reg}<16'b0110000111001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000111001000)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0110000111001001) && ({row_reg, col_reg}<16'b0110000111001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110000111001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110000111001100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110000111001101) && ({row_reg, col_reg}<16'b0110000111001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110000111001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110000111010000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110000111010001) && ({row_reg, col_reg}<16'b0110000111010100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110000111010100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110000111010101) && ({row_reg, col_reg}<16'b0110000111011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110000111011000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110000111011001) && ({row_reg, col_reg}<16'b0110000111011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110000111011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110000111011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110000111011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110000111011110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110000111011111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110000111100000) && ({row_reg, col_reg}<16'b0110000111101000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110000111101000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110000111101001) && ({row_reg, col_reg}<16'b0110000111101011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110000111101011) && ({row_reg, col_reg}<16'b0110000111101110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110000111101110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110000111101111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110000111110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110000111110001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110000111110010) && ({row_reg, col_reg}<16'b0110000111111001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110000111111001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110000111111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110000111111011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110000111111100) && ({row_reg, col_reg}<16'b0110000111111110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110000111111110)) color_data = 12'b010100110010;

		if(({row_reg, col_reg}==16'b0110000111111111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110001000000000) && ({row_reg, col_reg}<16'b0110001000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001000000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110001000000110) && ({row_reg, col_reg}<16'b0110001000001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110001000001000) && ({row_reg, col_reg}<16'b0110001000001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110001000001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001000001101) && ({row_reg, col_reg}<16'b0110001000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001000010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001000010001) && ({row_reg, col_reg}<16'b0110001001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110001001100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001001100100) && ({row_reg, col_reg}<16'b0110001001101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001001101000) && ({row_reg, col_reg}<16'b0110001001101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110001001101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001001101011) && ({row_reg, col_reg}<16'b0110001001101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110001001101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001001101110) && ({row_reg, col_reg}<16'b0110001001111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001001111001) && ({row_reg, col_reg}<16'b0110001001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110001001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001001111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110001001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110001001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001001111111) && ({row_reg, col_reg}<16'b0110001010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001010000010) && ({row_reg, col_reg}<16'b0110001010010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110001010010011) && ({row_reg, col_reg}<16'b0110001010010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001010010101) && ({row_reg, col_reg}<16'b0110001010011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001010011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001010011110) && ({row_reg, col_reg}<16'b0110001010100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001010100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001010100001) && ({row_reg, col_reg}<16'b0110001010100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110001010100011) && ({row_reg, col_reg}<16'b0110001010100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001010100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110001010100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001010100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110001010101000) && ({row_reg, col_reg}<16'b0110001010101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001010101011) && ({row_reg, col_reg}<16'b0110001010101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110001010101110) && ({row_reg, col_reg}<16'b0110001010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110001010110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110001010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001010110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110001010110110) && ({row_reg, col_reg}<16'b0110001010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110001010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110001010111001) && ({row_reg, col_reg}<16'b0110001010111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110001010111011) && ({row_reg, col_reg}<16'b0110001010111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110001010111101) && ({row_reg, col_reg}<16'b0110001011001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110001011001000) && ({row_reg, col_reg}<16'b0110001011001010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110001011001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001011001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001011001100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110001011001101) && ({row_reg, col_reg}<16'b0110001011001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110001011001111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110001011010000) && ({row_reg, col_reg}<16'b0110001011010101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110001011010101) && ({row_reg, col_reg}<16'b0110001011011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001011011000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110001011011001) && ({row_reg, col_reg}<16'b0110001011011011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110001011011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110001011011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110001011011101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110001011011110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110001011011111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110001011100000) && ({row_reg, col_reg}<16'b0110001011101001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110001011101001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110001011101010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110001011101011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110001011101100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110001011101101) && ({row_reg, col_reg}<16'b0110001011110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110001011110000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110001011110001) && ({row_reg, col_reg}<16'b0110001011111010)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110001011111010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110001011111011) && ({row_reg, col_reg}<16'b0110001011111110)) color_data = 12'b010101000011;

		if(({row_reg, col_reg}>=16'b0110001011111110) && ({row_reg, col_reg}<16'b0110001100000000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110001100000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001100000001) && ({row_reg, col_reg}<16'b0110001100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001100000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110001100000110) && ({row_reg, col_reg}<16'b0110001100001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110001100001000) && ({row_reg, col_reg}<16'b0110001100001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110001100001011) && ({row_reg, col_reg}<16'b0110001100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001100001101) && ({row_reg, col_reg}<16'b0110001100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110001100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001100010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001100010001) && ({row_reg, col_reg}<16'b0110001101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110001101100011) && ({row_reg, col_reg}<16'b0110001101101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001101101000) && ({row_reg, col_reg}<16'b0110001101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001101101011) && ({row_reg, col_reg}<16'b0110001101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110001101101101) && ({row_reg, col_reg}<16'b0110001101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001101111000) && ({row_reg, col_reg}<16'b0110001101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110001101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001101111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110001101111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110001101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001101111111) && ({row_reg, col_reg}<16'b0110001110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110001110000001) && ({row_reg, col_reg}<16'b0110001110010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110001110010011) && ({row_reg, col_reg}<16'b0110001110010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001110010101) && ({row_reg, col_reg}<16'b0110001110011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001110011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110001110011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001110011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001110100000) && ({row_reg, col_reg}<16'b0110001110100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110001110100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110001110100011) && ({row_reg, col_reg}<16'b0110001110100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110001110100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110001110100110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0110001110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110001110101000) && ({row_reg, col_reg}<16'b0110001110101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110001110101011) && ({row_reg, col_reg}<16'b0110001110101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110001110101110) && ({row_reg, col_reg}<16'b0110001110110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110001110110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110001110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001110110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110001110110110) && ({row_reg, col_reg}<16'b0110001110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110001110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110001110111001) && ({row_reg, col_reg}<16'b0110001110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001110111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110001110111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110001110111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110001110111110) && ({row_reg, col_reg}<16'b0110001111000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110001111000001) && ({row_reg, col_reg}<16'b0110001111000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110001111000100) && ({row_reg, col_reg}<16'b0110001111001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110001111001000)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==16'b0110001111001001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110001111001010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110001111001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001111001100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110001111001101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110001111001110) && ({row_reg, col_reg}<16'b0110001111010011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110001111010011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110001111010100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110001111010101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110001111010110) && ({row_reg, col_reg}<16'b0110001111011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110001111011101) && ({row_reg, col_reg}<16'b0110001111100000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110001111100000) && ({row_reg, col_reg}<16'b0110001111101001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110001111101001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110001111101010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110001111101011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110001111101100) && ({row_reg, col_reg}<16'b0110001111110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110001111110000) && ({row_reg, col_reg}<16'b0110001111110010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110001111110010) && ({row_reg, col_reg}<16'b0110001111110101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110001111110101) && ({row_reg, col_reg}<16'b0110001111111001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110001111111001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110001111111010) && ({row_reg, col_reg}<16'b0110001111111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110001111111100)) color_data = 12'b010101000010;

		if(({row_reg, col_reg}>=16'b0110001111111101) && ({row_reg, col_reg}<16'b0110010000000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110010000000000) && ({row_reg, col_reg}<16'b0110010000000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010000000010) && ({row_reg, col_reg}<16'b0110010000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010000000101) && ({row_reg, col_reg}<16'b0110010000000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110010000000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110010000001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110010000001001) && ({row_reg, col_reg}<16'b0110010000001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110010000001011) && ({row_reg, col_reg}<16'b0110010000001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110010000001101) && ({row_reg, col_reg}<16'b0110010000001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010000001111) && ({row_reg, col_reg}<16'b0110010000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010000010001) && ({row_reg, col_reg}<16'b0110010001100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110010001100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010001100011) && ({row_reg, col_reg}<16'b0110010001101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010001101001) && ({row_reg, col_reg}<16'b0110010001101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010001101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010001101101) && ({row_reg, col_reg}<16'b0110010001110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110010001110001) && ({row_reg, col_reg}<16'b0110010001110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010001110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010001110110) && ({row_reg, col_reg}<16'b0110010001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010001111000) && ({row_reg, col_reg}<16'b0110010001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010001111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110010001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110010001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110010001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010010000001) && ({row_reg, col_reg}<16'b0110010010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110010010010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010010010101) && ({row_reg, col_reg}<16'b0110010010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010010011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110010010100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110010010100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010010100010) && ({row_reg, col_reg}<16'b0110010010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010010100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010010100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110010010100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110010010100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110010010101000) && ({row_reg, col_reg}<16'b0110010010101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010010101011) && ({row_reg, col_reg}<16'b0110010010101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110010010101110) && ({row_reg, col_reg}<16'b0110010010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010010110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110010010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110010010110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110010010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110010010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010010110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110010010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110010010111001) && ({row_reg, col_reg}<16'b0110010010111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110010010111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110010010111100) && ({row_reg, col_reg}<16'b0110010010111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110010010111110) && ({row_reg, col_reg}<16'b0110010011000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110010011000010) && ({row_reg, col_reg}<16'b0110010011000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0110010011000100) && ({row_reg, col_reg}<16'b0110010011001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110010011001000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0110010011001001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110010011001010) && ({row_reg, col_reg}<16'b0110010011001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110010011001101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110010011001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110010011001111) && ({row_reg, col_reg}<16'b0110010011010011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110010011010011) && ({row_reg, col_reg}<16'b0110010011010110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110010011010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110010011010111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110010011011000) && ({row_reg, col_reg}<16'b0110010011011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110010011011010) && ({row_reg, col_reg}<16'b0110010011011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110010011011100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110010011011101) && ({row_reg, col_reg}<16'b0110010011100101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110010011100101) && ({row_reg, col_reg}<16'b0110010011100111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110010011100111) && ({row_reg, col_reg}<16'b0110010011101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110010011101001) && ({row_reg, col_reg}<16'b0110010011101011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110010011101011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110010011101100) && ({row_reg, col_reg}<16'b0110010011101111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110010011101111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110010011110000) && ({row_reg, col_reg}<16'b0110010011110010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110010011110010) && ({row_reg, col_reg}<16'b0110010011111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110010011111001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110010011111010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110010011111011) && ({row_reg, col_reg}<16'b0110010011111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110010011111101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110010011111110)) color_data = 12'b010000100001;

		if(({row_reg, col_reg}==16'b0110010011111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110010100000000) && ({row_reg, col_reg}<16'b0110010100000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110010100000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010100000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110010100000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010100000101) && ({row_reg, col_reg}<16'b0110010100000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110010100000111) && ({row_reg, col_reg}<16'b0110010100001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110010100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110010100001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110010100001011) && ({row_reg, col_reg}<16'b0110010100001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110010100001110) && ({row_reg, col_reg}<16'b0110010100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010100010001) && ({row_reg, col_reg}<16'b0110010101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110010101100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010101100011) && ({row_reg, col_reg}<16'b0110010101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010101101010) && ({row_reg, col_reg}<16'b0110010101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010101101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010101101101) && ({row_reg, col_reg}<16'b0110010101110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110010101110001) && ({row_reg, col_reg}<16'b0110010101111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110010101111001) && ({row_reg, col_reg}<16'b0110010101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010101111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110010101111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110010101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110010101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010110000001) && ({row_reg, col_reg}<16'b0110010110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110010110010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110010110010101) && ({row_reg, col_reg}<16'b0110010110011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010110011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110010110011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010110011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110010110011011) && ({row_reg, col_reg}<16'b0110010110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010110011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110010110100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110010110100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110010110100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010110100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110010110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010110100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110010110100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110010110100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110010110101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110010110101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110010110101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110010110101100) && ({row_reg, col_reg}<16'b0110010110101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110010110101110) && ({row_reg, col_reg}<16'b0110010110110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010110110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110010110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110010110110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110010110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110010110110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110010110110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110010110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110010110111001) && ({row_reg, col_reg}<16'b0110010110111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110010110111011) && ({row_reg, col_reg}<16'b0110010110111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110010110111111) && ({row_reg, col_reg}<16'b0110010111000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110010111000001) && ({row_reg, col_reg}<16'b0110010111000100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110010111000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0110010111000101) && ({row_reg, col_reg}<16'b0110010111001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110010111001000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0110010111001001) && ({row_reg, col_reg}<16'b0110010111001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110010111001011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110010111001100) && ({row_reg, col_reg}<16'b0110010111001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110010111001110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110010111001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110010111010000) && ({row_reg, col_reg}<16'b0110010111010011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110010111010011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110010111010100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110010111010101) && ({row_reg, col_reg}<16'b0110010111010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110010111010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110010111011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110010111011001) && ({row_reg, col_reg}<16'b0110010111100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110010111100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110010111100001) && ({row_reg, col_reg}<16'b0110010111101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110010111101100) && ({row_reg, col_reg}<16'b0110010111101110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110010111101110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110010111101111) && ({row_reg, col_reg}<16'b0110010111110100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110010111110100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110010111110101) && ({row_reg, col_reg}<16'b0110010111111011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110010111111011) && ({row_reg, col_reg}<16'b0110010111111101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110010111111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110010111111110)) color_data = 12'b010000100001;

		if(({row_reg, col_reg}==16'b0110010111111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011000000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011000000001) && ({row_reg, col_reg}<16'b0110011000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011000000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110011000000110) && ({row_reg, col_reg}<16'b0110011000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110011000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110011000001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110011000001011) && ({row_reg, col_reg}<16'b0110011000001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110011000001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011000001111) && ({row_reg, col_reg}<16'b0110011000010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110011000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011000010010) && ({row_reg, col_reg}<16'b0110011001100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110011001100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011001100011) && ({row_reg, col_reg}<16'b0110011001101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011001101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110011001101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011001101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110011001101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011001101110) && ({row_reg, col_reg}<16'b0110011001110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011001110010) && ({row_reg, col_reg}<16'b0110011001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011001111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110011001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110011001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110011001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011010000001) && ({row_reg, col_reg}<16'b0110011010010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110011010010101) && ({row_reg, col_reg}<16'b0110011010011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011010011000) && ({row_reg, col_reg}<16'b0110011010011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011010011010) && ({row_reg, col_reg}<16'b0110011010100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011010100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110011010100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110011010100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011010100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110011010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011010100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110011010100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110011010100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110011010101000) && ({row_reg, col_reg}<16'b0110011010101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110011010101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110011010101100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0110011010101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110011010101110) && ({row_reg, col_reg}<16'b0110011010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110011010110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110011010110011) && ({row_reg, col_reg}<16'b0110011010110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110011010110110) && ({row_reg, col_reg}<16'b0110011010111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110011010111000) && ({row_reg, col_reg}<16'b0110011010111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110011010111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110011010111100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0110011010111101) && ({row_reg, col_reg}<16'b0110011010111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110011010111111) && ({row_reg, col_reg}<16'b0110011011000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110011011000001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110011011000010) && ({row_reg, col_reg}<16'b0110011011000100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110011011000100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0110011011000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110011011000110) && ({row_reg, col_reg}<16'b0110011011001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110011011001000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011011001001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110011011001010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011011001011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110011011001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110011011001101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110011011001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110011011001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011011010000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110011011010001) && ({row_reg, col_reg}<16'b0110011011010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011011010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110011011011000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110011011011001) && ({row_reg, col_reg}<16'b0110011011011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110011011011011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110011011011100) && ({row_reg, col_reg}<16'b0110011011100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110011011100010) && ({row_reg, col_reg}<16'b0110011011100100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110011011100100) && ({row_reg, col_reg}<16'b0110011011100110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110011011100110) && ({row_reg, col_reg}<16'b0110011011101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110011011101001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110011011101010) && ({row_reg, col_reg}<16'b0110011011101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110011011101110) && ({row_reg, col_reg}<16'b0110011011110000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110011011110000) && ({row_reg, col_reg}<16'b0110011011110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011011110010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110011011110011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110011011110100) && ({row_reg, col_reg}<16'b0110011011111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110011011111001) && ({row_reg, col_reg}<16'b0110011011111011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110011011111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110011011111100) && ({row_reg, col_reg}<16'b0110011011111110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110011011111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0110011011111111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110011100000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011100000001) && ({row_reg, col_reg}<16'b0110011100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011100000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110011100000110) && ({row_reg, col_reg}<16'b0110011100001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110011100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110011100001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110011100001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011100001101) && ({row_reg, col_reg}<16'b0110011100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011100001111) && ({row_reg, col_reg}<16'b0110011100010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110011100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011100010010) && ({row_reg, col_reg}<16'b0110011101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110011101100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011101100011) && ({row_reg, col_reg}<16'b0110011101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011101101011) && ({row_reg, col_reg}<16'b0110011101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110011101101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110011101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011101101111) && ({row_reg, col_reg}<16'b0110011101110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011101110010) && ({row_reg, col_reg}<16'b0110011101110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011101110101) && ({row_reg, col_reg}<16'b0110011101110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011101110111) && ({row_reg, col_reg}<16'b0110011101111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011101111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110011101111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110011101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110011101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110011110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011110000001) && ({row_reg, col_reg}<16'b0110011110010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110011110010101) && ({row_reg, col_reg}<16'b0110011110011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110011110011001) && ({row_reg, col_reg}<16'b0110011110011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011110011011) && ({row_reg, col_reg}<16'b0110011110011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110011110011101) && ({row_reg, col_reg}<16'b0110011110100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110011110100000) && ({row_reg, col_reg}<16'b0110011110100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110011110100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110011110100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110011110100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110011110100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110011110100110) && ({row_reg, col_reg}<16'b0110011110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110011110101000) && ({row_reg, col_reg}<16'b0110011110101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110011110101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110011110101100) && ({row_reg, col_reg}<16'b0110011110101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110011110101110) && ({row_reg, col_reg}<16'b0110011110110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110011110110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110011110110011) && ({row_reg, col_reg}<16'b0110011110110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110011110110110) && ({row_reg, col_reg}<16'b0110011110111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110011110111000) && ({row_reg, col_reg}<16'b0110011110111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110011110111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110011110111100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0110011110111101) && ({row_reg, col_reg}<16'b0110011110111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110011110111111) && ({row_reg, col_reg}<16'b0110011111000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110011111000010) && ({row_reg, col_reg}<16'b0110011111000100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110011111000100) && ({row_reg, col_reg}<16'b0110011111000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110011111000111) && ({row_reg, col_reg}<16'b0110011111001001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110011111001001) && ({row_reg, col_reg}<16'b0110011111001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011111001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110011111001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110011111001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110011111001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110011111001111) && ({row_reg, col_reg}<16'b0110011111010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011111010001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110011111010010) && ({row_reg, col_reg}<16'b0110011111010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110011111010101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110011111010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011111010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110011111011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110011111011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110011111011010) && ({row_reg, col_reg}<16'b0110011111100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110011111100000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110011111100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110011111100010) && ({row_reg, col_reg}<16'b0110011111100100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110011111100100) && ({row_reg, col_reg}<16'b0110011111100110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110011111100110) && ({row_reg, col_reg}<16'b0110011111101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110011111101011) && ({row_reg, col_reg}<16'b0110011111110011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110011111110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110011111110100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110011111110101) && ({row_reg, col_reg}<16'b0110011111111111)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0110011111111111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110100000000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100000000001) && ({row_reg, col_reg}<16'b0110100000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100000000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110100000000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110100000000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110100000001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110100000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110100000001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110100000001011) && ({row_reg, col_reg}<16'b0110100000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100000001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110100000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100000010010) && ({row_reg, col_reg}<16'b0110100001100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110100001100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100001100011) && ({row_reg, col_reg}<16'b0110100001101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100001101001) && ({row_reg, col_reg}<16'b0110100001101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100001101011) && ({row_reg, col_reg}<16'b0110100001101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110100001101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110100001101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100001101111) && ({row_reg, col_reg}<16'b0110100001110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100001110011) && ({row_reg, col_reg}<16'b0110100001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100001111100) && ({row_reg, col_reg}<16'b0110100001111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110100001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110100001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100010000001) && ({row_reg, col_reg}<16'b0110100010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110100010010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100010010101) && ({row_reg, col_reg}<16'b0110100010011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110100010011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100010011010) && ({row_reg, col_reg}<16'b0110100010011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100010011101) && ({row_reg, col_reg}<16'b0110100010100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100010100001) && ({row_reg, col_reg}<16'b0110100010100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100010100011) && ({row_reg, col_reg}<16'b0110100010100110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110100010100110) && ({row_reg, col_reg}<16'b0110100010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110100010101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110100010101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100010101010) && ({row_reg, col_reg}<16'b0110100010101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110100010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100010101110) && ({row_reg, col_reg}<16'b0110100010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100010110000) && ({row_reg, col_reg}<16'b0110100010111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110100010111100) && ({row_reg, col_reg}<16'b0110100011001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110100011001001) && ({row_reg, col_reg}<16'b0110100011001011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110100011001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110100011001100) && ({row_reg, col_reg}<16'b0110100011001110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110100011001110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0110100011001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110100011010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110100011010001) && ({row_reg, col_reg}<16'b0110100011010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110100011010101) && ({row_reg, col_reg}<16'b0110100011010111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0110100011010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110100011011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110100011011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110100011011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110100011011011) && ({row_reg, col_reg}<16'b0110100011011101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110100011011101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110100011011110) && ({row_reg, col_reg}<16'b0110100011100000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110100011100000) && ({row_reg, col_reg}<16'b0110100011101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110100011101000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110100011101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110100011101010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110100011101011) && ({row_reg, col_reg}<16'b0110100011110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110100011110111) && ({row_reg, col_reg}<16'b0110100011111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110100011111011) && ({row_reg, col_reg}<16'b0110100011111110)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}>=16'b0110100011111110) && ({row_reg, col_reg}<16'b0110100100000000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110100100000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100100000001) && ({row_reg, col_reg}<16'b0110100100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100100000110) && ({row_reg, col_reg}<16'b0110100100001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110100100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110100100001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110100100001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100100001101) && ({row_reg, col_reg}<16'b0110100100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100100010010) && ({row_reg, col_reg}<16'b0110100101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110100101100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100101100011) && ({row_reg, col_reg}<16'b0110100101101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100101101000) && ({row_reg, col_reg}<16'b0110100101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100101101011) && ({row_reg, col_reg}<16'b0110100101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110100101101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100101101110) && ({row_reg, col_reg}<16'b0110100101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100101110000) && ({row_reg, col_reg}<16'b0110100101110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100101110100) && ({row_reg, col_reg}<16'b0110100101110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100101110111) && ({row_reg, col_reg}<16'b0110100101111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100101111001) && ({row_reg, col_reg}<16'b0110100101111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100101111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110100101111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110100101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110100101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100110000001) && ({row_reg, col_reg}<16'b0110100110010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110100110010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110100110010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100110010101) && ({row_reg, col_reg}<16'b0110100110011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110100110011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100110011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110100110011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110100110011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100110011101) && ({row_reg, col_reg}<16'b0110100110100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110100110100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110100110100001) && ({row_reg, col_reg}<16'b0110100110100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110100110100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110100110100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110100110100101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0110100110100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110100110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110100110101000) && ({row_reg, col_reg}<16'b0110100110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100110101011) && ({row_reg, col_reg}<16'b0110100110101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110100110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110100110101110) && ({row_reg, col_reg}<16'b0110100110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110100110110000) && ({row_reg, col_reg}<16'b0110100110110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110100110110010) && ({row_reg, col_reg}<16'b0110100111001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110100111001010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110100111001011) && ({row_reg, col_reg}<16'b0110100111001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110100111001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110100111001110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110100111001111) && ({row_reg, col_reg}<16'b0110100111010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110100111010010) && ({row_reg, col_reg}<16'b0110100111010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110100111010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110100111010101) && ({row_reg, col_reg}<16'b0110100111010111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110100111010111) && ({row_reg, col_reg}<16'b0110100111011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110100111011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110100111011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110100111011011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110100111011100) && ({row_reg, col_reg}<16'b0110100111011110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110100111011110) && ({row_reg, col_reg}<16'b0110100111100001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110100111100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110100111100010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110100111100011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110100111100100) && ({row_reg, col_reg}<16'b0110100111101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110100111101101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110100111101110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110100111101111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110100111110000) && ({row_reg, col_reg}<16'b0110100111110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110100111110110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110100111110111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110100111111000) && ({row_reg, col_reg}<16'b0110100111111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110100111111011) && ({row_reg, col_reg}<16'b0110100111111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110100111111101)) color_data = 12'b010100110010;

		if(({row_reg, col_reg}>=16'b0110100111111110) && ({row_reg, col_reg}<16'b0110101000000000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110101000000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101000000001) && ({row_reg, col_reg}<16'b0110101000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101000000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110101000000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110101000001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110101000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110101000001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110101000001011) && ({row_reg, col_reg}<16'b0110101000001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110101000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101000001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101000001111) && ({row_reg, col_reg}<16'b0110101000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101000010010) && ({row_reg, col_reg}<16'b0110101001100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110101001100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101001100011) && ({row_reg, col_reg}<16'b0110101001101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101001101000) && ({row_reg, col_reg}<16'b0110101001101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110101001101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101001101011) && ({row_reg, col_reg}<16'b0110101001101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101001101110) && ({row_reg, col_reg}<16'b0110101001110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101001110000) && ({row_reg, col_reg}<16'b0110101001110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110101001110100) && ({row_reg, col_reg}<16'b0110101001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101001111000) && ({row_reg, col_reg}<16'b0110101001111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110101001111010) && ({row_reg, col_reg}<16'b0110101001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101001111100) && ({row_reg, col_reg}<16'b0110101001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110101001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101010000001) && ({row_reg, col_reg}<16'b0110101010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110101010010100) && ({row_reg, col_reg}<16'b0110101010011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101010011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110101010011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101010011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110101010011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110101010011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101010011101) && ({row_reg, col_reg}<16'b0110101010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101010011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110101010100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110101010100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101010100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110101010100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110101010100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110101010100101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0110101010100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101010100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110101010101000) && ({row_reg, col_reg}<16'b0110101010101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110101010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101010101011) && ({row_reg, col_reg}<16'b0110101010101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110101010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101010101110) && ({row_reg, col_reg}<16'b0110101010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110101010110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110101010110001) && ({row_reg, col_reg}<16'b0110101010110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101010110011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110101010110100) && ({row_reg, col_reg}<16'b0110101010111101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110101010111101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110101010111110) && ({row_reg, col_reg}<16'b0110101011001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110101011001010) && ({row_reg, col_reg}<16'b0110101011001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110101011001101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110101011001110)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}>=16'b0110101011001111) && ({row_reg, col_reg}<16'b0110101011010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110101011010111) && ({row_reg, col_reg}<16'b0110101011011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110101011011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110101011011010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110101011011011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110101011011100) && ({row_reg, col_reg}<16'b0110101011011111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110101011011111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110101011100000) && ({row_reg, col_reg}<16'b0110101011100011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110101011100011) && ({row_reg, col_reg}<16'b0110101011100110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110101011100110) && ({row_reg, col_reg}<16'b0110101011101011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110101011101011) && ({row_reg, col_reg}<16'b0110101011101101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110101011101101) && ({row_reg, col_reg}<16'b0110101011110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110101011110000) && ({row_reg, col_reg}<16'b0110101011110110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110101011110110) && ({row_reg, col_reg}<16'b0110101011111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110101011111011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110101011111100) && ({row_reg, col_reg}<16'b0110101011111110)) color_data = 12'b010101000010;

		if(({row_reg, col_reg}>=16'b0110101011111110) && ({row_reg, col_reg}<16'b0110101100000000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110101100000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101100000001) && ({row_reg, col_reg}<16'b0110101100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101100000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110101100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110101100001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110101100001001) && ({row_reg, col_reg}<16'b0110101100001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110101100001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110101100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110101100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101100001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101100001111) && ({row_reg, col_reg}<16'b0110101100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101100010010) && ({row_reg, col_reg}<16'b0110101101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110101101100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101101100011) && ({row_reg, col_reg}<16'b0110101101100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101101100110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101101100111) && ({row_reg, col_reg}<16'b0110101101101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101101101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110101101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101101101011) && ({row_reg, col_reg}<16'b0110101101101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110101101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101101101111) && ({row_reg, col_reg}<16'b0110101101110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110101101110011) && ({row_reg, col_reg}<16'b0110101101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101101111000) && ({row_reg, col_reg}<16'b0110101101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110101101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101101111100) && ({row_reg, col_reg}<16'b0110101101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101101111110) && ({row_reg, col_reg}<16'b0110101110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101110000001) && ({row_reg, col_reg}<16'b0110101110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110101110010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101110010101) && ({row_reg, col_reg}<16'b0110101110011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110101110011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110101110011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110101110011100) && ({row_reg, col_reg}<16'b0110101110011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110101110011110) && ({row_reg, col_reg}<16'b0110101110100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110101110100000) && ({row_reg, col_reg}<16'b0110101110100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110101110100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110101110100011) && ({row_reg, col_reg}<16'b0110101110100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110101110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110101110100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110101110101000) && ({row_reg, col_reg}<16'b0110101110101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110101110101011) && ({row_reg, col_reg}<16'b0110101110101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110101110101110) && ({row_reg, col_reg}<16'b0110101110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110101110110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110101110110001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0110101110110010) && ({row_reg, col_reg}<16'b0110101110110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110101110110100) && ({row_reg, col_reg}<16'b0110101110111000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110101110111000) && ({row_reg, col_reg}<16'b0110101110111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110101110111110) && ({row_reg, col_reg}<16'b0110101111000001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110101111000001) && ({row_reg, col_reg}<16'b0110101111000100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110101111000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110101111000101) && ({row_reg, col_reg}<16'b0110101111000111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110101111000111) && ({row_reg, col_reg}<16'b0110101111001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110101111001101) && ({row_reg, col_reg}<16'b0110101111001111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110101111001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110101111010000) && ({row_reg, col_reg}<16'b0110101111010100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110101111010100) && ({row_reg, col_reg}<16'b0110101111010110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110101111010110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110101111010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0110101111011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110101111011001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0110101111011010) && ({row_reg, col_reg}<16'b0110101111011100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110101111011100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110101111011101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110101111011110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110101111011111) && ({row_reg, col_reg}<16'b0110101111100010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110101111100010) && ({row_reg, col_reg}<16'b0110101111100101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110101111100101) && ({row_reg, col_reg}<16'b0110101111100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110101111100111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110101111101000) && ({row_reg, col_reg}<16'b0110101111101010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110101111101010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110101111101011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110101111101100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110101111101101) && ({row_reg, col_reg}<16'b0110101111110000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110101111110000) && ({row_reg, col_reg}<16'b0110101111110100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110101111110100) && ({row_reg, col_reg}<16'b0110101111110110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110101111110110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110101111110111) && ({row_reg, col_reg}<16'b0110101111111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110101111111100)) color_data = 12'b010100110010;

		if(({row_reg, col_reg}>=16'b0110101111111101) && ({row_reg, col_reg}<16'b0110110000000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110110000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110110000000001) && ({row_reg, col_reg}<16'b0110110000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110000000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110110000000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110110000001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110110000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110110000001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110110000001011) && ({row_reg, col_reg}<16'b0110110000001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110110000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110000001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110000001111) && ({row_reg, col_reg}<16'b0110110000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110000010010) && ({row_reg, col_reg}<16'b0110110001100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110001100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110001100011) && ({row_reg, col_reg}<16'b0110110001100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110001100110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110001100111) && ({row_reg, col_reg}<16'b0110110001101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110001101001) && ({row_reg, col_reg}<16'b0110110001101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110001101011) && ({row_reg, col_reg}<16'b0110110001101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110001101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110110001101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110001101111) && ({row_reg, col_reg}<16'b0110110001110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110001110001) && ({row_reg, col_reg}<16'b0110110001110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110001110111) && ({row_reg, col_reg}<16'b0110110001111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110001111010) && ({row_reg, col_reg}<16'b0110110001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110001111100) && ({row_reg, col_reg}<16'b0110110001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110001111110) && ({row_reg, col_reg}<16'b0110110010000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110110010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110010000001) && ({row_reg, col_reg}<16'b0110110010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110010010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110010010101) && ({row_reg, col_reg}<16'b0110110010011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110010011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110110010011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110110010011100) && ({row_reg, col_reg}<16'b0110110010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110010011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110110010100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110010100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110110010100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110110010100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110110010100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110110010100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110110010100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110010100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110110010101000) && ({row_reg, col_reg}<16'b0110110010101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110110010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110010101011) && ({row_reg, col_reg}<16'b0110110010101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110110010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110010101110) && ({row_reg, col_reg}<16'b0110110010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110110010110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110110010110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110110010110010) && ({row_reg, col_reg}<16'b0110110010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110110010110101) && ({row_reg, col_reg}<16'b0110110010111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110110010111010) && ({row_reg, col_reg}<16'b0110110011000001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110110011000001) && ({row_reg, col_reg}<16'b0110110011001000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110110011001000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110110011001001) && ({row_reg, col_reg}<16'b0110110011001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110011001101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110110011001110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0110110011001111) && ({row_reg, col_reg}<16'b0110110011010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110110011010101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110110011010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110110011010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110011011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110110011011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110110011011010) && ({row_reg, col_reg}<16'b0110110011011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110110011011100) && ({row_reg, col_reg}<16'b0110110011100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110110011100010) && ({row_reg, col_reg}<16'b0110110011100100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110110011100100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110110011100101) && ({row_reg, col_reg}<16'b0110110011100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0110110011100111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110110011101000) && ({row_reg, col_reg}<16'b0110110011101011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110110011101011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110110011101100) && ({row_reg, col_reg}<16'b0110110011101110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110110011101110) && ({row_reg, col_reg}<16'b0110110011110000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110110011110000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110110011110001) && ({row_reg, col_reg}<16'b0110110011110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110110011110011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110110011110100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110110011110101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0110110011110110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==16'b0110110011110111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110110011111000) && ({row_reg, col_reg}<16'b0110110011111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110110011111110)) color_data = 12'b010000100001;

		if(({row_reg, col_reg}==16'b0110110011111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110110100000001) && ({row_reg, col_reg}<16'b0110110100000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110100000011) && ({row_reg, col_reg}<16'b0110110100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110100000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110110100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110110100001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110110100001001) && ({row_reg, col_reg}<16'b0110110100001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110110100001011) && ({row_reg, col_reg}<16'b0110110100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110100001101) && ({row_reg, col_reg}<16'b0110110100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110100010010) && ({row_reg, col_reg}<16'b0110110101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110101100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110101100011) && ({row_reg, col_reg}<16'b0110110101101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110101101001) && ({row_reg, col_reg}<16'b0110110101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110101101011) && ({row_reg, col_reg}<16'b0110110101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110101101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110110101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110101110000) && ({row_reg, col_reg}<16'b0110110101111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110101111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110101111010) && ({row_reg, col_reg}<16'b0110110101111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110101111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110110101111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110101111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110110101111111) && ({row_reg, col_reg}<16'b0110110110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110110000001) && ({row_reg, col_reg}<16'b0110110110010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110110010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110110010100) && ({row_reg, col_reg}<16'b0110110110011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110110110011001) && ({row_reg, col_reg}<16'b0110110110011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110110110011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110110011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110110110011101) && ({row_reg, col_reg}<16'b0110110110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110110011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110110110100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110110110100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110110110100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110110110100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110110110100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110110110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110110110100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110110100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110110110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110110110101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110110110101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110110110101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110110110101100) && ({row_reg, col_reg}<16'b0110110110101110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110110110101110) && ({row_reg, col_reg}<16'b0110110110110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110110110110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110110110110001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0110110110110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110110110110011) && ({row_reg, col_reg}<16'b0110110110110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0110110110110111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0110110110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110110110111001) && ({row_reg, col_reg}<16'b0110110111000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110111000000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110110111000001) && ({row_reg, col_reg}<16'b0110110111001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110110111001001) && ({row_reg, col_reg}<16'b0110110111001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110110111001100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110110111001101) && ({row_reg, col_reg}<16'b0110110111001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110111001111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0110110111010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110110111010001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0110110111010010) && ({row_reg, col_reg}<16'b0110110111010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110110111010100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110110111010101) && ({row_reg, col_reg}<16'b0110110111010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110110111010111) && ({row_reg, col_reg}<16'b0110110111011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110110111011111) && ({row_reg, col_reg}<16'b0110110111100001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110110111100001) && ({row_reg, col_reg}<16'b0110110111100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110110111100011) && ({row_reg, col_reg}<16'b0110110111100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110110111100101) && ({row_reg, col_reg}<16'b0110110111100111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0110110111100111) && ({row_reg, col_reg}<16'b0110110111101010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110110111101010) && ({row_reg, col_reg}<16'b0110110111101101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110110111101101) && ({row_reg, col_reg}<16'b0110110111101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110110111101111) && ({row_reg, col_reg}<16'b0110110111110001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110110111110001) && ({row_reg, col_reg}<16'b0110110111110011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110110111110011) && ({row_reg, col_reg}<16'b0110110111110101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0110110111110101) && ({row_reg, col_reg}<16'b0110110111111000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110110111111000) && ({row_reg, col_reg}<16'b0110110111111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110110111111011)) color_data = 12'b010000110001;

		if(({row_reg, col_reg}>=16'b0110110111111100) && ({row_reg, col_reg}<16'b0110111000000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110111000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110111000000001) && ({row_reg, col_reg}<16'b0110111000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111000000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110111000000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0110111000001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110111000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110111000001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110111000001011) && ({row_reg, col_reg}<16'b0110111000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111000010010) && ({row_reg, col_reg}<16'b0110111001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110111001100011) && ({row_reg, col_reg}<16'b0110111001101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111001101000) && ({row_reg, col_reg}<16'b0110111001101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111001101011) && ({row_reg, col_reg}<16'b0110111001101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110111001101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110111001101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111001101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111001110000) && ({row_reg, col_reg}<16'b0110111001111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111001111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111001111010) && ({row_reg, col_reg}<16'b0110111001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111001111100) && ({row_reg, col_reg}<16'b0110111001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111001111110) && ({row_reg, col_reg}<16'b0110111010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111010000010) && ({row_reg, col_reg}<16'b0110111010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110111010010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111010010101) && ({row_reg, col_reg}<16'b0110111010011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111010011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110111010011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110111010011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111010011101) && ({row_reg, col_reg}<16'b0110111010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111010011111) && ({row_reg, col_reg}<16'b0110111010100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110111010100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111010100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110111010100011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0110111010100100) && ({row_reg, col_reg}<16'b0110111010100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111010100110) && ({row_reg, col_reg}<16'b0110111010101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110111010101000) && ({row_reg, col_reg}<16'b0110111010101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111010101011) && ({row_reg, col_reg}<16'b0110111010101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110111010101101) && ({row_reg, col_reg}<16'b0110111010110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110111010110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110111010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111010110100) && ({row_reg, col_reg}<16'b0110111010111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110111010111001) && ({row_reg, col_reg}<16'b0110111010111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111010111100) && ({row_reg, col_reg}<16'b0110111011000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110111011000001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110111011000010) && ({row_reg, col_reg}<16'b0110111011001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110111011001101) && ({row_reg, col_reg}<16'b0110111011011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110111011011010) && ({row_reg, col_reg}<16'b0110111011011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111011011100) && ({row_reg, col_reg}<16'b0110111011100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110111011100010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110111011100011) && ({row_reg, col_reg}<16'b0110111011101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110111011101001) && ({row_reg, col_reg}<16'b0110111011110100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110111011110100) && ({row_reg, col_reg}<16'b0110111011111000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111011111000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110111011111001) && ({row_reg, col_reg}<16'b0110111011111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110111011111101)) color_data = 12'b001000100001;

		if(({row_reg, col_reg}>=16'b0110111011111110) && ({row_reg, col_reg}<16'b0110111100000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110111100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110111100000001) && ({row_reg, col_reg}<16'b0110111100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111100000110) && ({row_reg, col_reg}<16'b0110111100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111100001010) && ({row_reg, col_reg}<16'b0110111100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111100010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111100010001) && ({row_reg, col_reg}<16'b0110111101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110111101100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111101100100) && ({row_reg, col_reg}<16'b0110111101101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111101101000) && ({row_reg, col_reg}<16'b0110111101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110111101101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110111101101101) && ({row_reg, col_reg}<16'b0110111101101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111101110000) && ({row_reg, col_reg}<16'b0110111101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0110111101111000) && ({row_reg, col_reg}<16'b0110111101111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111101111010) && ({row_reg, col_reg}<16'b0110111110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111110000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111110000010) && ({row_reg, col_reg}<16'b0110111110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110111110010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111110010101) && ({row_reg, col_reg}<16'b0110111110011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111110011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0110111110011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110111110011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0110111110011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0110111110011101) && ({row_reg, col_reg}<16'b0110111110100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111110100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0110111110100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0110111110100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0110111110100011) && ({row_reg, col_reg}<16'b0110111110100101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0110111110100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111110100110) && ({row_reg, col_reg}<16'b0110111110101110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110111110101110) && ({row_reg, col_reg}<16'b0110111110110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0110111110110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110111110110011) && ({row_reg, col_reg}<16'b0110111110110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111110110110) && ({row_reg, col_reg}<16'b0110111110111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0110111110111100) && ({row_reg, col_reg}<16'b0110111110111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0110111110111111) && ({row_reg, col_reg}<16'b0110111111000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0110111111000010) && ({row_reg, col_reg}<16'b0110111111001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0110111111001101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110111111001110) && ({row_reg, col_reg}<16'b0110111111100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110111111100111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110111111101000) && ({row_reg, col_reg}<16'b0110111111101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110111111101100) && ({row_reg, col_reg}<16'b0110111111101111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0110111111101111) && ({row_reg, col_reg}<16'b0110111111110100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0110111111110100) && ({row_reg, col_reg}<16'b0110111111110110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0110111111110110) && ({row_reg, col_reg}<16'b0110111111111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0110111111111101)) color_data = 12'b001000100001;

		if(({row_reg, col_reg}>=16'b0110111111111110) && ({row_reg, col_reg}<16'b0111000000000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111000000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000000000001) && ({row_reg, col_reg}<16'b0111000000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000000000110) && ({row_reg, col_reg}<16'b0111000000001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000000001011) && ({row_reg, col_reg}<16'b0111000000001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111000000001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111000000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000000010000) && ({row_reg, col_reg}<16'b0111000000010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111000000010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000000010100) && ({row_reg, col_reg}<16'b0111000001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111000001100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000001100100) && ({row_reg, col_reg}<16'b0111000001101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000001101001) && ({row_reg, col_reg}<16'b0111000001101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111000001101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000001101101) && ({row_reg, col_reg}<16'b0111000001101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111000001101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000001110000) && ({row_reg, col_reg}<16'b0111000001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000001111000) && ({row_reg, col_reg}<16'b0111000001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000001111011) && ({row_reg, col_reg}<16'b0111000010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000010000001) && ({row_reg, col_reg}<16'b0111000010010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000010010101) && ({row_reg, col_reg}<16'b0111000010011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000010011000) && ({row_reg, col_reg}<16'b0111000010011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111000010011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111000010011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000010011100) && ({row_reg, col_reg}<16'b0111000010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111000010100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000010100100) && ({row_reg, col_reg}<16'b0111000010100110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111000010100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000010100111) && ({row_reg, col_reg}<16'b0111000010101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111000010101101) && ({row_reg, col_reg}<16'b0111000010101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111000010101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111000010110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000010110001) && ({row_reg, col_reg}<16'b0111000010110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111000010110110) && ({row_reg, col_reg}<16'b0111000010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111000010111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111000010111001) && ({row_reg, col_reg}<16'b0111000010111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111000010111100) && ({row_reg, col_reg}<16'b0111000010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111000010111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111000010111111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0111000011000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000011000001) && ({row_reg, col_reg}<16'b0111000011000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111000011000100) && ({row_reg, col_reg}<16'b0111000011001101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111000011001101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111000011001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111000011001111) && ({row_reg, col_reg}<16'b0111000011010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000011010001) && ({row_reg, col_reg}<16'b0111000011010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111000011010011) && ({row_reg, col_reg}<16'b0111000011010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111000011010110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111000011010111) && ({row_reg, col_reg}<16'b0111000011011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111000011011010) && ({row_reg, col_reg}<16'b0111000011011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111000011011101) && ({row_reg, col_reg}<16'b0111000011100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111000011100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000011100110) && ({row_reg, col_reg}<16'b0111000011101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111000011101011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111000011101100) && ({row_reg, col_reg}<16'b0111000011110000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111000011110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111000011110001)) color_data = 12'b010000100001;

		if(({row_reg, col_reg}>=16'b0111000011110010) && ({row_reg, col_reg}<16'b0111000100000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111000100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111000100000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000100000010) && ({row_reg, col_reg}<16'b0111000100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000100000101) && ({row_reg, col_reg}<16'b0111000100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000100001011) && ({row_reg, col_reg}<16'b0111000100001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111000100001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111000100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000100010000) && ({row_reg, col_reg}<16'b0111000100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111000100010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000100010100) && ({row_reg, col_reg}<16'b0111000101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111000101100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000101100011) && ({row_reg, col_reg}<16'b0111000101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111000101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000101101011) && ({row_reg, col_reg}<16'b0111000101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111000101101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111000101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111000101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000101110000) && ({row_reg, col_reg}<16'b0111000101111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000101111001) && ({row_reg, col_reg}<16'b0111000101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000101111011) && ({row_reg, col_reg}<16'b0111000110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111000110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000110000001) && ({row_reg, col_reg}<16'b0111000110010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111000110010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000110010110) && ({row_reg, col_reg}<16'b0111000110011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111000110011010) && ({row_reg, col_reg}<16'b0111000110011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111000110011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000110011101) && ({row_reg, col_reg}<16'b0111000110100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111000110100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111000110100001) && ({row_reg, col_reg}<16'b0111000110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111000110100100) && ({row_reg, col_reg}<16'b0111000110101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111000110101000) && ({row_reg, col_reg}<16'b0111000110101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111000110101011) && ({row_reg, col_reg}<16'b0111000110110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000110110000) && ({row_reg, col_reg}<16'b0111000110110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111000110110110) && ({row_reg, col_reg}<16'b0111000110111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111000110111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111000110111010) && ({row_reg, col_reg}<16'b0111000110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000110111110) && ({row_reg, col_reg}<16'b0111000111000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111000111000000) && ({row_reg, col_reg}<16'b0111000111000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000111000010) && ({row_reg, col_reg}<16'b0111000111000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111000111000110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111000111000111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111000111001000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111000111001001) && ({row_reg, col_reg}<16'b0111000111001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111000111001100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111000111001101) && ({row_reg, col_reg}<16'b0111000111001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111000111001111) && ({row_reg, col_reg}<16'b0111000111010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000111010001) && ({row_reg, col_reg}<16'b0111000111010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111000111010011) && ({row_reg, col_reg}<16'b0111000111011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111000111011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111000111011111) && ({row_reg, col_reg}<16'b0111000111100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111000111100110) && ({row_reg, col_reg}<16'b0111000111101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111000111101000) && ({row_reg, col_reg}<16'b0111000111111100)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}>=16'b0111000111111100) && ({row_reg, col_reg}<16'b0111001000000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001000000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001000000010) && ({row_reg, col_reg}<16'b0111001000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001000000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001000000111) && ({row_reg, col_reg}<16'b0111001000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111001000001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001000001010) && ({row_reg, col_reg}<16'b0111001000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001000010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001000010001) && ({row_reg, col_reg}<16'b0111001001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111001001100011) && ({row_reg, col_reg}<16'b0111001001101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001001101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001001101011) && ({row_reg, col_reg}<16'b0111001001101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001001101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111001001101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001001101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001001110000) && ({row_reg, col_reg}<16'b0111001001111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001001111001) && ({row_reg, col_reg}<16'b0111001001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001001111011) && ({row_reg, col_reg}<16'b0111001001111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001001111110) && ({row_reg, col_reg}<16'b0111001010000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001010000001) && ({row_reg, col_reg}<16'b0111001010010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111001010010101) && ({row_reg, col_reg}<16'b0111001010010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001010010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001010011000) && ({row_reg, col_reg}<16'b0111001010011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001010011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001010011100) && ({row_reg, col_reg}<16'b0111001010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001010100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111001010100101) && ({row_reg, col_reg}<16'b0111001010101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001010101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111001010101001) && ({row_reg, col_reg}<16'b0111001010101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001010101100) && ({row_reg, col_reg}<16'b0111001010101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0111001010101110) && ({row_reg, col_reg}<16'b0111001010110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111001010110110) && ({row_reg, col_reg}<16'b0111001010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001010111000) && ({row_reg, col_reg}<16'b0111001010111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001010111101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001010111110) && ({row_reg, col_reg}<16'b0111001011000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111001011000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111001011000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111001011000010) && ({row_reg, col_reg}<16'b0111001011000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111001011000100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0111001011000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001011000110) && ({row_reg, col_reg}<16'b0111001011001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111001011001010) && ({row_reg, col_reg}<16'b0111001011001100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111001011001100) && ({row_reg, col_reg}<16'b0111001011001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111001011001110) && ({row_reg, col_reg}<16'b0111001011010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111001011010000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0111001011010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111001011010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001011010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001011010100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111001011010101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111001011010110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111001011010111) && ({row_reg, col_reg}<16'b0111001011011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001011011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111001011011111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111001011100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001011100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111001011100010) && ({row_reg, col_reg}<16'b0111001011100100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111001011100100) && ({row_reg, col_reg}<16'b0111001011110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001011110111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111001011111000) && ({row_reg, col_reg}<16'b0111001011111011)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}>=16'b0111001011111011) && ({row_reg, col_reg}<16'b0111001100000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001100000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001100000010) && ({row_reg, col_reg}<16'b0111001100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001100000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111001100000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001100001000) && ({row_reg, col_reg}<16'b0111001100001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111001100001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111001100001011) && ({row_reg, col_reg}<16'b0111001100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001100010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001100010001) && ({row_reg, col_reg}<16'b0111001101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111001101100011) && ({row_reg, col_reg}<16'b0111001101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001101101011) && ({row_reg, col_reg}<16'b0111001101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001101101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111001101101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001101101111) && ({row_reg, col_reg}<16'b0111001101110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001101110001) && ({row_reg, col_reg}<16'b0111001101111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001101111001) && ({row_reg, col_reg}<16'b0111001101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111001101111011) && ({row_reg, col_reg}<16'b0111001110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001110000001) && ({row_reg, col_reg}<16'b0111001110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111001110010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111001110010101) && ({row_reg, col_reg}<16'b0111001110011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001110011110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111001110011111) && ({row_reg, col_reg}<16'b0111001110100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111001110100010) && ({row_reg, col_reg}<16'b0111001110100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111001110100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111001110100101) && ({row_reg, col_reg}<16'b0111001110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111001110101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111001110101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111001110101100) && ({row_reg, col_reg}<16'b0111001110101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001110101110) && ({row_reg, col_reg}<16'b0111001110110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111001110110110) && ({row_reg, col_reg}<16'b0111001110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001110111000) && ({row_reg, col_reg}<16'b0111001110111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001110111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001111000000) && ({row_reg, col_reg}<16'b0111001111000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111001111000011) && ({row_reg, col_reg}<16'b0111001111000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111001111000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001111001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001111001001) && ({row_reg, col_reg}<16'b0111001111001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111001111001110) && ({row_reg, col_reg}<16'b0111001111010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111001111010001) && ({row_reg, col_reg}<16'b0111001111010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001111010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001111010100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111001111010101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=16'b0111001111010110) && ({row_reg, col_reg}<16'b0111001111011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001111011000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111001111011001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111001111011010) && ({row_reg, col_reg}<16'b0111001111011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001111011110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111001111011111) && ({row_reg, col_reg}<16'b0111001111100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001111100001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111001111100010) && ({row_reg, col_reg}<16'b0111001111100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111001111100111) && ({row_reg, col_reg}<16'b0111001111101010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111001111101010) && ({row_reg, col_reg}<16'b0111001111110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111001111110010) && ({row_reg, col_reg}<16'b0111001111110110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111001111110110) && ({row_reg, col_reg}<16'b0111001111111000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111001111111000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111001111111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111001111111010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111001111111011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111001111111100) && ({row_reg, col_reg}<16'b0111001111111111)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0111001111111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111010000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111010000000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010000000010) && ({row_reg, col_reg}<16'b0111010000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010000000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111010000000111) && ({row_reg, col_reg}<16'b0111010000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111010000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111010000001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111010000001011) && ({row_reg, col_reg}<16'b0111010000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010000010001) && ({row_reg, col_reg}<16'b0111010001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111010001100011) && ({row_reg, col_reg}<16'b0111010001101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010001101001) && ({row_reg, col_reg}<16'b0111010001101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111010001101011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==16'b0111010001101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111010001101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010001101110) && ({row_reg, col_reg}<16'b0111010010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010010000001) && ({row_reg, col_reg}<16'b0111010010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111010010010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010010010101) && ({row_reg, col_reg}<16'b0111010010010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010010010111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111010010011000) && ({row_reg, col_reg}<16'b0111010010011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111010010011010) && ({row_reg, col_reg}<16'b0111010010100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010010100000) && ({row_reg, col_reg}<16'b0111010010100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111010010100110) && ({row_reg, col_reg}<16'b0111010010101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010010101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111010010101101) && ({row_reg, col_reg}<16'b0111010010101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111010010101111) && ({row_reg, col_reg}<16'b0111010011000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111010011000100) && ({row_reg, col_reg}<16'b0111010011001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111010011001010) && ({row_reg, col_reg}<16'b0111010011001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111010011001100) && ({row_reg, col_reg}<16'b0111010011001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111010011001111) && ({row_reg, col_reg}<16'b0111010011010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111010011010010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0111010011010011) && ({row_reg, col_reg}<16'b0111010011010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111010011010101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==16'b0111010011010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111010011010111) && ({row_reg, col_reg}<16'b0111010011011001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111010011011001) && ({row_reg, col_reg}<16'b0111010011011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111010011011111) && ({row_reg, col_reg}<16'b0111010011100001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111010011100001) && ({row_reg, col_reg}<16'b0111010011101011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111010011101011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111010011101100) && ({row_reg, col_reg}<16'b0111010011110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111010011110001) && ({row_reg, col_reg}<16'b0111010011111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111010011111001) && ({row_reg, col_reg}<16'b0111010011111100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111010011111100) && ({row_reg, col_reg}<16'b0111010011111111)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0111010011111111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111010100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111010100000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010100000010) && ({row_reg, col_reg}<16'b0111010100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010100000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111010100000111) && ({row_reg, col_reg}<16'b0111010100001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111010100001010) && ({row_reg, col_reg}<16'b0111010100001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010100001100) && ({row_reg, col_reg}<16'b0111010100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111010100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010100010010) && ({row_reg, col_reg}<16'b0111010101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111010101100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010101100100) && ({row_reg, col_reg}<16'b0111010101101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010101101001) && ({row_reg, col_reg}<16'b0111010101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111010101101100) && ({row_reg, col_reg}<16'b0111010110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111010110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010110000001) && ({row_reg, col_reg}<16'b0111010110010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111010110010011) && ({row_reg, col_reg}<16'b0111010110010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111010110010101) && ({row_reg, col_reg}<16'b0111010110011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010110011000) && ({row_reg, col_reg}<16'b0111010110011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111010110011010) && ({row_reg, col_reg}<16'b0111010110101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111010110101000) && ({row_reg, col_reg}<16'b0111010110101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111010110101100) && ({row_reg, col_reg}<16'b0111010110101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111010110101111) && ({row_reg, col_reg}<16'b0111010110110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111010110110001) && ({row_reg, col_reg}<16'b0111010111000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111010111000110) && ({row_reg, col_reg}<16'b0111010111001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111010111001010) && ({row_reg, col_reg}<16'b0111010111001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111010111001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111010111001101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0111010111001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111010111001111) && ({row_reg, col_reg}<16'b0111010111010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111010111010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111010111010011)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0111010111010100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111010111010101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111010111010110) && ({row_reg, col_reg}<16'b0111010111100011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111010111100011) && ({row_reg, col_reg}<16'b0111010111100101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111010111100101) && ({row_reg, col_reg}<16'b0111010111101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111010111101100) && ({row_reg, col_reg}<16'b0111010111101110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111010111101110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111010111101111) && ({row_reg, col_reg}<16'b0111010111110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111010111110010) && ({row_reg, col_reg}<16'b0111010111110100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111010111110100) && ({row_reg, col_reg}<16'b0111010111111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111010111111010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111010111111011)) color_data = 12'b010000110001;

		if(({row_reg, col_reg}>=16'b0111010111111100) && ({row_reg, col_reg}<16'b0111011000000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111011000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111011000000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011000000010) && ({row_reg, col_reg}<16'b0111011000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011000000110) && ({row_reg, col_reg}<16'b0111011000001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011000001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111011000001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011000001010) && ({row_reg, col_reg}<16'b0111011000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011000001110) && ({row_reg, col_reg}<16'b0111011000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011000010010) && ({row_reg, col_reg}<16'b0111011001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111011001100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111011001100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011001100101) && ({row_reg, col_reg}<16'b0111011001101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111011001101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011001101001) && ({row_reg, col_reg}<16'b0111011001101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011001101011) && ({row_reg, col_reg}<16'b0111011001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011001111000) && ({row_reg, col_reg}<16'b0111011001111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011001111010) && ({row_reg, col_reg}<16'b0111011001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011001111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011010000001) && ({row_reg, col_reg}<16'b0111011010010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111011010010010) && ({row_reg, col_reg}<16'b0111011010010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011010010100) && ({row_reg, col_reg}<16'b0111011010011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011010011000) && ({row_reg, col_reg}<16'b0111011010011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011010011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111011010011100) && ({row_reg, col_reg}<16'b0111011010011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111011010011110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111011010011111) && ({row_reg, col_reg}<16'b0111011010100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011010100010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111011010100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111011010100100) && ({row_reg, col_reg}<16'b0111011010101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111011010101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011010101011) && ({row_reg, col_reg}<16'b0111011010110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111011010110001) && ({row_reg, col_reg}<16'b0111011010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111011010110011) && ({row_reg, col_reg}<16'b0111011010110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111011010110110) && ({row_reg, col_reg}<16'b0111011010111000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111011010111000) && ({row_reg, col_reg}<16'b0111011011001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111011011001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111011011001101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0111011011001110) && ({row_reg, col_reg}<16'b0111011011010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111011011010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0111011011010011) && ({row_reg, col_reg}<16'b0111011011010110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}>=16'b0111011011010110) && ({row_reg, col_reg}<16'b0111011011101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111011011101100) && ({row_reg, col_reg}<16'b0111011011101110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111011011101110) && ({row_reg, col_reg}<16'b0111011011110001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111011011110001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111011011110010) && ({row_reg, col_reg}<16'b0111011011110100)) color_data = 12'b010101000010;

		if(({row_reg, col_reg}>=16'b0111011011110100) && ({row_reg, col_reg}<16'b0111011100000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111011100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111011100000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011100000010) && ({row_reg, col_reg}<16'b0111011100000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011100000111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111011100001000) && ({row_reg, col_reg}<16'b0111011100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011100001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011100001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011100001110) && ({row_reg, col_reg}<16'b0111011100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011100010001) && ({row_reg, col_reg}<16'b0111011101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111011101100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011101100100) && ({row_reg, col_reg}<16'b0111011101101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011101101000) && ({row_reg, col_reg}<16'b0111011101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011101101011) && ({row_reg, col_reg}<16'b0111011101110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011101110111) && ({row_reg, col_reg}<16'b0111011101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011101111011) && ({row_reg, col_reg}<16'b0111011101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011101111111) && ({row_reg, col_reg}<16'b0111011110000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011110000010) && ({row_reg, col_reg}<16'b0111011110000100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011110000100) && ({row_reg, col_reg}<16'b0111011110001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011110001000) && ({row_reg, col_reg}<16'b0111011110001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011110001100) && ({row_reg, col_reg}<16'b0111011110001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011110001110) && ({row_reg, col_reg}<16'b0111011110010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011110010010) && ({row_reg, col_reg}<16'b0111011110011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111011110011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111011110011001) && ({row_reg, col_reg}<16'b0111011110011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011110011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111011110011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111011110011110)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b0111011110011111) && ({row_reg, col_reg}<16'b0111011110100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011110100010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111011110100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111011110100100) && ({row_reg, col_reg}<16'b0111011110100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111011110100111) && ({row_reg, col_reg}<16'b0111011110101001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111011110101001) && ({row_reg, col_reg}<16'b0111011110101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111011110101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111011110101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111011110101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111011110101110) && ({row_reg, col_reg}<16'b0111011110110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111011110110000) && ({row_reg, col_reg}<16'b0111011110110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111011110110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111011110110100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111011110110101) && ({row_reg, col_reg}<16'b0111011111001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111011111001110) && ({row_reg, col_reg}<16'b0111011111010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111011111010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111011111010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111011111010011) && ({row_reg, col_reg}<16'b0111011111010110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111011111010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111011111010111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111011111011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111011111011001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111011111011010) && ({row_reg, col_reg}<16'b0111011111101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111011111101100) && ({row_reg, col_reg}<16'b0111011111101110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111011111101110) && ({row_reg, col_reg}<16'b0111011111110010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111011111110010) && ({row_reg, col_reg}<16'b0111011111110101)) color_data = 12'b010100110010;

		if(({row_reg, col_reg}>=16'b0111011111110101) && ({row_reg, col_reg}<16'b0111100000000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111100000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111100000000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111100000000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111100000000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111100000000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111100000000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100000000110) && ({row_reg, col_reg}<16'b0111100000001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111100000001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111100000001001) && ({row_reg, col_reg}<16'b0111100000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100000001100) && ({row_reg, col_reg}<16'b0111100000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100000001111) && ({row_reg, col_reg}<16'b0111100000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100000010001) && ({row_reg, col_reg}<16'b0111100001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111100001100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111100001100100) && ({row_reg, col_reg}<16'b0111100001100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100001100110) && ({row_reg, col_reg}<16'b0111100001101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100001101011) && ({row_reg, col_reg}<16'b0111100001101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111100001101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100001110000) && ({row_reg, col_reg}<16'b0111100001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100001111000) && ({row_reg, col_reg}<16'b0111100001111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100001111010) && ({row_reg, col_reg}<16'b0111100010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100010000000) && ({row_reg, col_reg}<16'b0111100010000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100010000010) && ({row_reg, col_reg}<16'b0111100010010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100010010111) && ({row_reg, col_reg}<16'b0111100010011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111100010011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100010011011) && ({row_reg, col_reg}<16'b0111100010100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111100010100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111100010100111) && ({row_reg, col_reg}<16'b0111100010101001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111100010101001) && ({row_reg, col_reg}<16'b0111100010101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100010101011) && ({row_reg, col_reg}<16'b0111100010101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111100010101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111100010101110) && ({row_reg, col_reg}<16'b0111100010110001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111100010110001) && ({row_reg, col_reg}<16'b0111100010110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100010110011) && ({row_reg, col_reg}<16'b0111100010110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111100010110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111100010110110) && ({row_reg, col_reg}<16'b0111100011000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111100011000000) && ({row_reg, col_reg}<16'b0111100011000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111100011000010) && ({row_reg, col_reg}<16'b0111100011001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111100011001111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0111100011010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111100011010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111100011010010)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==16'b0111100011010011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==16'b0111100011010100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==16'b0111100011010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111100011010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b0111100011010111) && ({row_reg, col_reg}<16'b0111100011011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111100011011001) && ({row_reg, col_reg}<16'b0111100011011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111100011011011)) color_data = 12'b010000100001;

		if(({row_reg, col_reg}>=16'b0111100011011100) && ({row_reg, col_reg}<16'b0111100100000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111100100000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111100100000001) && ({row_reg, col_reg}<16'b0111100100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111100100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100100000110) && ({row_reg, col_reg}<16'b0111100100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111100100001001) && ({row_reg, col_reg}<16'b0111100100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100100001101) && ({row_reg, col_reg}<16'b0111100100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111100100010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111100100010001) && ({row_reg, col_reg}<16'b0111100100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111100100100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111100100100100) && ({row_reg, col_reg}<16'b0111100101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111100101100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111100101100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100101100100) && ({row_reg, col_reg}<16'b0111100101100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111100101100110) && ({row_reg, col_reg}<16'b0111100101101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111100101101000) && ({row_reg, col_reg}<16'b0111100101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100101101010) && ({row_reg, col_reg}<16'b0111100101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100101101100) && ({row_reg, col_reg}<16'b0111100101111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100101111001) && ({row_reg, col_reg}<16'b0111100101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100101111011) && ({row_reg, col_reg}<16'b0111100101111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111100101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111100101111111) && ({row_reg, col_reg}<16'b0111100110010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100110010100) && ({row_reg, col_reg}<16'b0111100110010111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111100110010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100110011000) && ({row_reg, col_reg}<16'b0111100110011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111100110011011) && ({row_reg, col_reg}<16'b0111100110011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100110011101) && ({row_reg, col_reg}<16'b0111100110100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100110100101) && ({row_reg, col_reg}<16'b0111100110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111100110101000) && ({row_reg, col_reg}<16'b0111100110101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100110101011) && ({row_reg, col_reg}<16'b0111100110101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b0111100110101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111100110101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111100110101111) && ({row_reg, col_reg}<16'b0111100110110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111100110110001) && ({row_reg, col_reg}<16'b0111100110110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111100110110100) && ({row_reg, col_reg}<16'b0111100110110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111100110110111) && ({row_reg, col_reg}<16'b0111100110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111100110111010) && ({row_reg, col_reg}<16'b0111100110111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111100110111111) && ({row_reg, col_reg}<16'b0111100111000011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111100111000011) && ({row_reg, col_reg}<16'b0111100111001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111100111001101)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=16'b0111100111001110) && ({row_reg, col_reg}<16'b0111100111010010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111100111010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111100111010011)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111100111010100) && ({row_reg, col_reg}<16'b0111100111010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111100111010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111100111010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111100111011000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111100111011001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0111100111011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111100111011011) && ({row_reg, col_reg}<16'b0111100111011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111100111011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111100111100000) && ({row_reg, col_reg}<16'b0111100111111001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111100111111001)) color_data = 12'b010100110010;

		if(({row_reg, col_reg}>=16'b0111100111111010) && ({row_reg, col_reg}<16'b0111101000000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111101000000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101000000001) && ({row_reg, col_reg}<16'b0111101000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101000000101) && ({row_reg, col_reg}<16'b0111101000000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101000000111) && ({row_reg, col_reg}<16'b0111101000001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111101000001010) && ({row_reg, col_reg}<16'b0111101000001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111101000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101000001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111101000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101000010000) && ({row_reg, col_reg}<16'b0111101000100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101000100101) && ({row_reg, col_reg}<16'b0111101001010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111101001010010) && ({row_reg, col_reg}<16'b0111101001100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111101001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111101001100010) && ({row_reg, col_reg}<16'b0111101001100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101001100100) && ({row_reg, col_reg}<16'b0111101001101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111101001101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101001101010) && ({row_reg, col_reg}<16'b0111101001101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101001101101) && ({row_reg, col_reg}<16'b0111101001110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101001110100) && ({row_reg, col_reg}<16'b0111101001110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101001110110) && ({row_reg, col_reg}<16'b0111101001111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111101001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101001111001) && ({row_reg, col_reg}<16'b0111101001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101001111011) && ({row_reg, col_reg}<16'b0111101001111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101001111111) && ({row_reg, col_reg}<16'b0111101010010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101010010100) && ({row_reg, col_reg}<16'b0111101010010111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101010010111) && ({row_reg, col_reg}<16'b0111101010011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101010011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101010011100) && ({row_reg, col_reg}<16'b0111101010011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101010011110) && ({row_reg, col_reg}<16'b0111101010100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101010100101) && ({row_reg, col_reg}<16'b0111101010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111101010101000) && ({row_reg, col_reg}<16'b0111101010101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111101010101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111101010101100) && ({row_reg, col_reg}<16'b0111101010101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0111101010101110) && ({row_reg, col_reg}<16'b0111101010110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111101010110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101010110010) && ({row_reg, col_reg}<16'b0111101010110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111101010110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101010110110) && ({row_reg, col_reg}<16'b0111101010111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111101010111011) && ({row_reg, col_reg}<16'b0111101010111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101010111111) && ({row_reg, col_reg}<16'b0111101011000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111101011000010) && ({row_reg, col_reg}<16'b0111101011001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101011001000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111101011001001) && ({row_reg, col_reg}<16'b0111101011001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101011001101) && ({row_reg, col_reg}<16'b0111101011010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111101011010001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0111101011010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101011010011) && ({row_reg, col_reg}<16'b0111101011010101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111101011010101) && ({row_reg, col_reg}<16'b0111101011010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101011010111) && ({row_reg, col_reg}<16'b0111101011011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111101011011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101011100000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111101011100001) && ({row_reg, col_reg}<16'b0111101011111111)) color_data = 12'b010000110010;

		if(({row_reg, col_reg}==16'b0111101011111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111101100000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101100000001) && ({row_reg, col_reg}<16'b0111101100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101100000101) && ({row_reg, col_reg}<16'b0111101100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111101100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111101100001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111101100001011) && ({row_reg, col_reg}<16'b0111101100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101100001101) && ({row_reg, col_reg}<16'b0111101100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101100001111) && ({row_reg, col_reg}<16'b0111101100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101100010001) && ({row_reg, col_reg}<16'b0111101100010110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111101100010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111101100010111) && ({row_reg, col_reg}<16'b0111101100100100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101100100100) && ({row_reg, col_reg}<16'b0111101101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111101101010011) && ({row_reg, col_reg}<16'b0111101101010111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111101101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111101101011000) && ({row_reg, col_reg}<16'b0111101101011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111101101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111101101011100) && ({row_reg, col_reg}<16'b0111101101100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101101100010) && ({row_reg, col_reg}<16'b0111101101100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101101100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111101101100101) && ({row_reg, col_reg}<16'b0111101101100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111101101100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111101101101000) && ({row_reg, col_reg}<16'b0111101101101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101101101100) && ({row_reg, col_reg}<16'b0111101101110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101101110101) && ({row_reg, col_reg}<16'b0111101101110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101101110111) && ({row_reg, col_reg}<16'b0111101101111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101101111111) && ({row_reg, col_reg}<16'b0111101110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101110000001) && ({row_reg, col_reg}<16'b0111101110001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101110001000) && ({row_reg, col_reg}<16'b0111101110001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101110001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111101110001011) && ({row_reg, col_reg}<16'b0111101110011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101110011100) && ({row_reg, col_reg}<16'b0111101110011110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111101110011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111101110011111) && ({row_reg, col_reg}<16'b0111101110100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101110100010) && ({row_reg, col_reg}<16'b0111101110101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111101110101011) && ({row_reg, col_reg}<16'b0111101110110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111101110110001) && ({row_reg, col_reg}<16'b0111101110110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101110110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111101110111000) && ({row_reg, col_reg}<16'b0111101110111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111101110111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111101110111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111101110111101) && ({row_reg, col_reg}<16'b0111101110111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101110111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111101111000000) && ({row_reg, col_reg}<16'b0111101111000010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111101111000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111101111000011) && ({row_reg, col_reg}<16'b0111101111000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101111000111) && ({row_reg, col_reg}<16'b0111101111001001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111101111001001) && ({row_reg, col_reg}<16'b0111101111001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101111001100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111101111001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101111001110) && ({row_reg, col_reg}<16'b0111101111010001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b0111101111010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101111010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111101111010011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111101111010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111101111010101) && ({row_reg, col_reg}<16'b0111101111011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111101111011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111101111011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101111011010) && ({row_reg, col_reg}<16'b0111101111011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111101111011100) && ({row_reg, col_reg}<16'b0111101111011110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0111101111011110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111101111011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111101111100000) && ({row_reg, col_reg}<16'b0111101111100100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101111100100) && ({row_reg, col_reg}<16'b0111101111100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111101111100111) && ({row_reg, col_reg}<16'b0111101111101001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=16'b0111101111101001) && ({row_reg, col_reg}<16'b0111101111101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111101111101100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111101111101101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111101111101110) && ({row_reg, col_reg}<16'b0111101111110010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111101111110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111101111110011) && ({row_reg, col_reg}<16'b0111101111110110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111101111110110) && ({row_reg, col_reg}<16'b0111101111111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111101111111011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111101111111100)) color_data = 12'b010000100001;

		if(({row_reg, col_reg}>=16'b0111101111111101) && ({row_reg, col_reg}<16'b0111110000000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111110000000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110000000001) && ({row_reg, col_reg}<16'b0111110000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110000000110) && ({row_reg, col_reg}<16'b0111110000001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110000001001) && ({row_reg, col_reg}<16'b0111110000001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111110000001011) && ({row_reg, col_reg}<16'b0111110000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110000001101) && ({row_reg, col_reg}<16'b0111110000001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110000001111) && ({row_reg, col_reg}<16'b0111110000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110000010001) && ({row_reg, col_reg}<16'b0111110000010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110000010101) && ({row_reg, col_reg}<16'b0111110000011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111110000011000) && ({row_reg, col_reg}<16'b0111110000100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110000100011) && ({row_reg, col_reg}<16'b0111110001010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111110001010100) && ({row_reg, col_reg}<16'b0111110001010110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110001010110) && ({row_reg, col_reg}<16'b0111110001011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111110001011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110001011110) && ({row_reg, col_reg}<16'b0111110001100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111110001100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111110001100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110001100100) && ({row_reg, col_reg}<16'b0111110001100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110001100110) && ({row_reg, col_reg}<16'b0111110001110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110001110110) && ({row_reg, col_reg}<16'b0111110001111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110001111000) && ({row_reg, col_reg}<16'b0111110001111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111110001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110010000000) && ({row_reg, col_reg}<16'b0111110010001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110010001000) && ({row_reg, col_reg}<16'b0111110010011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110010011101) && ({row_reg, col_reg}<16'b0111110010011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110010011111) && ({row_reg, col_reg}<16'b0111110010100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110010100010) && ({row_reg, col_reg}<16'b0111110010100100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111110010100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111110010100101) && ({row_reg, col_reg}<16'b0111110010101011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111110010101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110010101100) && ({row_reg, col_reg}<16'b0111110010101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110010101110) && ({row_reg, col_reg}<16'b0111110010110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111110010110000) && ({row_reg, col_reg}<16'b0111110010111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111110010111000) && ({row_reg, col_reg}<16'b0111110010111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110010111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111110010111101) && ({row_reg, col_reg}<16'b0111110010111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110010111111) && ({row_reg, col_reg}<16'b0111110011000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110011000111) && ({row_reg, col_reg}<16'b0111110011001001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111110011001001) && ({row_reg, col_reg}<16'b0111110011001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111110011001111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b0111110011010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110011010001) && ({row_reg, col_reg}<16'b0111110011010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111110011010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111110011010100) && ({row_reg, col_reg}<16'b0111110011011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110011011011) && ({row_reg, col_reg}<16'b0111110011011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111110011011110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111110011011111) && ({row_reg, col_reg}<16'b0111110011100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111110011100001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0111110011100010) && ({row_reg, col_reg}<16'b0111110011100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110011100100) && ({row_reg, col_reg}<16'b0111110011100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110011100111) && ({row_reg, col_reg}<16'b0111110011101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111110011101100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111110011101101) && ({row_reg, col_reg}<16'b0111110011110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111110011110000) && ({row_reg, col_reg}<16'b0111110011110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110011110011) && ({row_reg, col_reg}<16'b0111110011110110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111110011110110) && ({row_reg, col_reg}<16'b0111110011111000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111110011111000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111110011111001) && ({row_reg, col_reg}<16'b0111110011111110)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}>=16'b0111110011111110) && ({row_reg, col_reg}<16'b0111110100000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111110100000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110100000001) && ({row_reg, col_reg}<16'b0111110100000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110100000011) && ({row_reg, col_reg}<16'b0111110100000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111110100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110100000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111110100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0111110100001000) && ({row_reg, col_reg}<16'b0111110100001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111110100001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111110100001011) && ({row_reg, col_reg}<16'b0111110100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110100010001) && ({row_reg, col_reg}<16'b0111110100010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110100010100) && ({row_reg, col_reg}<16'b0111110101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111110101100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110101100100) && ({row_reg, col_reg}<16'b0111110101100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110101100110) && ({row_reg, col_reg}<16'b0111110101101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111110101101000) && ({row_reg, col_reg}<16'b0111110101101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110101101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110101101101) && ({row_reg, col_reg}<16'b0111110101110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110101110111) && ({row_reg, col_reg}<16'b0111110101111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110101111001) && ({row_reg, col_reg}<16'b0111110110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110110000000) && ({row_reg, col_reg}<16'b0111110110000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110110000010) && ({row_reg, col_reg}<16'b0111110110000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110110000111) && ({row_reg, col_reg}<16'b0111110110001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111110110001010) && ({row_reg, col_reg}<16'b0111110110011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110110011110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111110110011111) && ({row_reg, col_reg}<16'b0111110110100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111110110100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111110110100100) && ({row_reg, col_reg}<16'b0111110110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110110101000) && ({row_reg, col_reg}<16'b0111110110101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111110110101010) && ({row_reg, col_reg}<16'b0111110110101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111110110101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110110101101) && ({row_reg, col_reg}<16'b0111110110101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111110110101111) && ({row_reg, col_reg}<16'b0111110110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110110110011) && ({row_reg, col_reg}<16'b0111110110110110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0111110110110110) && ({row_reg, col_reg}<16'b0111110110111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111110110111001) && ({row_reg, col_reg}<16'b0111110110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111110110111101) && ({row_reg, col_reg}<16'b0111110110111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111110110111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110111000000) && ({row_reg, col_reg}<16'b0111110111000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111110111000111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111110111001000) && ({row_reg, col_reg}<16'b0111110111010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111110111010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111110111010011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b0111110111010100) && ({row_reg, col_reg}<16'b0111110111010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111110111010111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111110111011000) && ({row_reg, col_reg}<16'b0111110111011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110111011011) && ({row_reg, col_reg}<16'b0111110111011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110111011101) && ({row_reg, col_reg}<16'b0111110111011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110111011111) && ({row_reg, col_reg}<16'b0111110111100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110111100100) && ({row_reg, col_reg}<16'b0111110111100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111110111100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111110111100111) && ({row_reg, col_reg}<16'b0111110111101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111110111101010) && ({row_reg, col_reg}<16'b0111110111101100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111110111101100) && ({row_reg, col_reg}<16'b0111110111101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111110111101110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111110111101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111110111110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111110111110001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111110111110010) && ({row_reg, col_reg}<16'b0111110111110111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111110111110111) && ({row_reg, col_reg}<16'b0111110111111001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111110111111001) && ({row_reg, col_reg}<16'b0111110111111011)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}>=16'b0111110111111011) && ({row_reg, col_reg}<16'b0111111000000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111000000000) && ({row_reg, col_reg}<16'b0111111000000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111000000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111111000000111) && ({row_reg, col_reg}<16'b0111111000001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111111000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111111000001010) && ({row_reg, col_reg}<16'b0111111000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111000010001) && ({row_reg, col_reg}<16'b0111111000010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111111000010100) && ({row_reg, col_reg}<16'b0111111001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111111001100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111001100100) && ({row_reg, col_reg}<16'b0111111001110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111001110111) && ({row_reg, col_reg}<16'b0111111001111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111001111001) && ({row_reg, col_reg}<16'b0111111010001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111010001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111010001010) && ({row_reg, col_reg}<16'b0111111010011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111010011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111111010011001) && ({row_reg, col_reg}<16'b0111111010011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111010011110) && ({row_reg, col_reg}<16'b0111111010100001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111111010100001) && ({row_reg, col_reg}<16'b0111111010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111010100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111111010100101) && ({row_reg, col_reg}<16'b0111111010101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111111010101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111111010101001) && ({row_reg, col_reg}<16'b0111111010101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111010101100) && ({row_reg, col_reg}<16'b0111111010101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111111010101111) && ({row_reg, col_reg}<16'b0111111010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111010111000) && ({row_reg, col_reg}<16'b0111111010111011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111111010111011) && ({row_reg, col_reg}<16'b0111111011000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111111011000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111111011000100) && ({row_reg, col_reg}<16'b0111111011000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111011000110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111111011000111) && ({row_reg, col_reg}<16'b0111111011010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111011010000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b0111111011010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111011010010) && ({row_reg, col_reg}<16'b0111111011010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111111011010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111111011010101) && ({row_reg, col_reg}<16'b0111111011010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111011010111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111111011011000) && ({row_reg, col_reg}<16'b0111111011011010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111111011011010) && ({row_reg, col_reg}<16'b0111111011100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111011100000) && ({row_reg, col_reg}<16'b0111111011100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111011100100) && ({row_reg, col_reg}<16'b0111111011101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111111011101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111011101001) && ({row_reg, col_reg}<16'b0111111011101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111011101101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b0111111011101110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b0111111011101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111011110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111111011110001) && ({row_reg, col_reg}<16'b0111111011110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b0111111011110110) && ({row_reg, col_reg}<16'b0111111011111001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111011111001) && ({row_reg, col_reg}<16'b0111111011111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111111011111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111111011111100) && ({row_reg, col_reg}<16'b0111111011111110)) color_data = 12'b001000100001;

		if(({row_reg, col_reg}>=16'b0111111011111110) && ({row_reg, col_reg}<16'b0111111100000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111100000000) && ({row_reg, col_reg}<16'b0111111100000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111111100000010) && ({row_reg, col_reg}<16'b0111111100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111100000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111111100000111) && ({row_reg, col_reg}<16'b0111111100001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111100001001) && ({row_reg, col_reg}<16'b0111111100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111111100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111100001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b0111111100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111100010000) && ({row_reg, col_reg}<16'b0111111100010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111111100010100) && ({row_reg, col_reg}<16'b0111111101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b0111111101100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111101100100) && ({row_reg, col_reg}<16'b0111111101110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111101110111) && ({row_reg, col_reg}<16'b0111111101111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111101111001) && ({row_reg, col_reg}<16'b0111111101111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111101111100) && ({row_reg, col_reg}<16'b0111111101111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111111101111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111101111111) && ({row_reg, col_reg}<16'b0111111110000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b0111111110000010) && ({row_reg, col_reg}<16'b0111111110000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111110000101) && ({row_reg, col_reg}<16'b0111111110000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111110000111) && ({row_reg, col_reg}<16'b0111111110001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111110001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111110001100) && ({row_reg, col_reg}<16'b0111111110010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111110010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111110010001) && ({row_reg, col_reg}<16'b0111111110010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111110010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b0111111110010110) && ({row_reg, col_reg}<16'b0111111110100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111110100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b0111111110100110) && ({row_reg, col_reg}<16'b0111111110101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111111110101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0111111110101001) && ({row_reg, col_reg}<16'b0111111110110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b0111111110110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111111110110001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b0111111110110010) && ({row_reg, col_reg}<16'b0111111110110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111110110110) && ({row_reg, col_reg}<16'b0111111110111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111111110111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b0111111110111010) && ({row_reg, col_reg}<16'b0111111110111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b0111111110111101) && ({row_reg, col_reg}<16'b0111111110111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111111110111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b0111111111000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111111111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111111000010) && ({row_reg, col_reg}<16'b0111111111000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111111111000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111111000101) && ({row_reg, col_reg}<16'b0111111111001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111111001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111111111001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111111010000) && ({row_reg, col_reg}<16'b0111111111010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111111111010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b0111111111010011) && ({row_reg, col_reg}<16'b0111111111010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b0111111111010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b0111111111010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111111010111) && ({row_reg, col_reg}<16'b0111111111011010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111111111011010) && ({row_reg, col_reg}<16'b0111111111100100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111111100100) && ({row_reg, col_reg}<16'b0111111111101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111111101001) && ({row_reg, col_reg}<16'b0111111111110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b0111111111110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b0111111111110001) && ({row_reg, col_reg}<16'b0111111111110100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b0111111111110100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b0111111111110101) && ({row_reg, col_reg}<16'b0111111111110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b0111111111110111) && ({row_reg, col_reg}<16'b0111111111111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b0111111111111001) && ({row_reg, col_reg}<16'b0111111111111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b0111111111111011)) color_data = 12'b001000010001;

		if(({row_reg, col_reg}>=16'b0111111111111100) && ({row_reg, col_reg}<16'b1000000000000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000000000000) && ({row_reg, col_reg}<16'b1000000000000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000000000000010) && ({row_reg, col_reg}<16'b1000000000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000000000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000000000000111) && ({row_reg, col_reg}<16'b1000000000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000000000001001) && ({row_reg, col_reg}<16'b1000000000001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000000000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000000001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000000000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000000010000) && ({row_reg, col_reg}<16'b1000000000010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000000000010011) && ({row_reg, col_reg}<16'b1000000001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000000001100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000000001100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000001100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000000001100110) && ({row_reg, col_reg}<16'b1000000001101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000001101011) && ({row_reg, col_reg}<16'b1000000001101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000001101101) && ({row_reg, col_reg}<16'b1000000001110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000001110111) && ({row_reg, col_reg}<16'b1000000001111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000001111001) && ({row_reg, col_reg}<16'b1000000001111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000000001111111) && ({row_reg, col_reg}<16'b1000000010000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000000010000010) && ({row_reg, col_reg}<16'b1000000010000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000010000101) && ({row_reg, col_reg}<16'b1000000010000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000010000111) && ({row_reg, col_reg}<16'b1000000010001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000010001010) && ({row_reg, col_reg}<16'b1000000010001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000010001100) && ({row_reg, col_reg}<16'b1000000010001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000010001111) && ({row_reg, col_reg}<16'b1000000010010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000010010001) && ({row_reg, col_reg}<16'b1000000010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000010100100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000000010100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000010100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000000010100111) && ({row_reg, col_reg}<16'b1000000010101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000010101011) && ({row_reg, col_reg}<16'b1000000010101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000000010101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000000010101110)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b1000000010101111) && ({row_reg, col_reg}<16'b1000000010110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000000010110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000010110010) && ({row_reg, col_reg}<16'b1000000010110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000010110110) && ({row_reg, col_reg}<16'b1000000010111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000010111000) && ({row_reg, col_reg}<16'b1000000010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000010111010) && ({row_reg, col_reg}<16'b1000000010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000000010111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000000010111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000000010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000010111111) && ({row_reg, col_reg}<16'b1000000011000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000000011000001) && ({row_reg, col_reg}<16'b1000000011000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000011000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000000011000101) && ({row_reg, col_reg}<16'b1000000011001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000011001001) && ({row_reg, col_reg}<16'b1000000011010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000000011010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000000011010011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000000011010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000011010101) && ({row_reg, col_reg}<16'b1000000011011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000011011000) && ({row_reg, col_reg}<16'b1000000011011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000000011011100) && ({row_reg, col_reg}<16'b1000000011100100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000011100100) && ({row_reg, col_reg}<16'b1000000011100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000000011100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000011100111) && ({row_reg, col_reg}<16'b1000000011101110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000011101110) && ({row_reg, col_reg}<16'b1000000011110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000000011110010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000000011110011) && ({row_reg, col_reg}<16'b1000000011110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000000011110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000011110111) && ({row_reg, col_reg}<16'b1000000011111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000000011111001) && ({row_reg, col_reg}<16'b1000000011111100)) color_data = 12'b001000100001;

		if(({row_reg, col_reg}>=16'b1000000011111100) && ({row_reg, col_reg}<16'b1000000100000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000000100000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000000100000001) && ({row_reg, col_reg}<16'b1000000100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000100000110) && ({row_reg, col_reg}<16'b1000000100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000000100001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000000100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000000100001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000100001011) && ({row_reg, col_reg}<16'b1000000100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000100001101) && ({row_reg, col_reg}<16'b1000000100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000100010001) && ({row_reg, col_reg}<16'b1000000100010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000000100010011) && ({row_reg, col_reg}<16'b1000000101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000000101100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000101100100) && ({row_reg, col_reg}<16'b1000000101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000101101010) && ({row_reg, col_reg}<16'b1000000101101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000101101101) && ({row_reg, col_reg}<16'b1000000101110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000101110111) && ({row_reg, col_reg}<16'b1000000101111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000101111001) && ({row_reg, col_reg}<16'b1000000101111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000101111100) && ({row_reg, col_reg}<16'b1000000101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000000101111110) && ({row_reg, col_reg}<16'b1000000110000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000000110000010) && ({row_reg, col_reg}<16'b1000000110010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000110010100) && ({row_reg, col_reg}<16'b1000000110011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000110011000) && ({row_reg, col_reg}<16'b1000000110100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000110100001) && ({row_reg, col_reg}<16'b1000000110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000110100100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000000110100101) && ({row_reg, col_reg}<16'b1000000110100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000000110100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000000110101000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000000110101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000000110101010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1000000110101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000000110101100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000000110101101) && ({row_reg, col_reg}<16'b1000000110101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000000110101111) && ({row_reg, col_reg}<16'b1000000110110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000110110001) && ({row_reg, col_reg}<16'b1000000110110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000110110011) && ({row_reg, col_reg}<16'b1000000110110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000110110110) && ({row_reg, col_reg}<16'b1000000110111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000000110111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000000110111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000000110111010) && ({row_reg, col_reg}<16'b1000000110111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000000110111100) && ({row_reg, col_reg}<16'b1000000110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000000110111111) && ({row_reg, col_reg}<16'b1000000111000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000000111000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000000111000100) && ({row_reg, col_reg}<16'b1000000111001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000000111001001) && ({row_reg, col_reg}<16'b1000000111001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000111001011) && ({row_reg, col_reg}<16'b1000000111011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000000111011000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000000111011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000111011010) && ({row_reg, col_reg}<16'b1000000111011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000000111011100) && ({row_reg, col_reg}<16'b1000000111101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000000111101100) && ({row_reg, col_reg}<16'b1000000111110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000111110001) && ({row_reg, col_reg}<16'b1000000111110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000000111110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000111110110) && ({row_reg, col_reg}<16'b1000000111111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000000111111000) && ({row_reg, col_reg}<16'b1000000111111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000000111111010) && ({row_reg, col_reg}<16'b1000000111111111)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}==16'b1000000111111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000001000000000) && ({row_reg, col_reg}<16'b1000001000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001000000110) && ({row_reg, col_reg}<16'b1000001000001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000001000001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001000001011) && ({row_reg, col_reg}<16'b1000001000001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001000001101) && ({row_reg, col_reg}<16'b1000001000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001000010001) && ({row_reg, col_reg}<16'b1000001000010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000001000010100) && ({row_reg, col_reg}<16'b1000001001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000001001100011) && ({row_reg, col_reg}<16'b1000001001100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000001001100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001001100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001001100111) && ({row_reg, col_reg}<16'b1000001001101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001001101010) && ({row_reg, col_reg}<16'b1000001001101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001001101101) && ({row_reg, col_reg}<16'b1000001001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001001111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001001111001) && ({row_reg, col_reg}<16'b1000001001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001001111100) && ({row_reg, col_reg}<16'b1000001010000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000001010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000001010000001) && ({row_reg, col_reg}<16'b1000001010000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001010000101) && ({row_reg, col_reg}<16'b1000001010000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001010000111) && ({row_reg, col_reg}<16'b1000001010010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001010010101) && ({row_reg, col_reg}<16'b1000001010010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001010010111) && ({row_reg, col_reg}<16'b1000001010011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001010011101) && ({row_reg, col_reg}<16'b1000001010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001010011111) && ({row_reg, col_reg}<16'b1000001010100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001010100010) && ({row_reg, col_reg}<16'b1000001010101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001010101001) && ({row_reg, col_reg}<16'b1000001010101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000001010101011) && ({row_reg, col_reg}<16'b1000001010101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000001010101110) && ({row_reg, col_reg}<16'b1000001010110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000001010110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001010110011) && ({row_reg, col_reg}<16'b1000001010110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001010110110) && ({row_reg, col_reg}<16'b1000001010111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000001010111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000001010111011)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=16'b1000001010111100) && ({row_reg, col_reg}<16'b1000001010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001010111110) && ({row_reg, col_reg}<16'b1000001011000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000001011000001) && ({row_reg, col_reg}<16'b1000001011000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000001011000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001011000101) && ({row_reg, col_reg}<16'b1000001011001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000001011001011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001011001100) && ({row_reg, col_reg}<16'b1000001011010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000001011010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000001011010011) && ({row_reg, col_reg}<16'b1000001011011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000001011011011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000001011011100) && ({row_reg, col_reg}<16'b1000001011101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001011101101) && ({row_reg, col_reg}<16'b1000001011110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001011110001) && ({row_reg, col_reg}<16'b1000001011110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000001011110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000001011110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001011110101) && ({row_reg, col_reg}<16'b1000001011111011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001011111011) && ({row_reg, col_reg}<16'b1000001011111110)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}>=16'b1000001011111110) && ({row_reg, col_reg}<16'b1000001100000000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000001100000000) && ({row_reg, col_reg}<16'b1000001100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001100000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000001100000111) && ({row_reg, col_reg}<16'b1000001100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000001100001001) && ({row_reg, col_reg}<16'b1000001100001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000001100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001100001101) && ({row_reg, col_reg}<16'b1000001100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001100010001) && ({row_reg, col_reg}<16'b1000001100010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000001100010100) && ({row_reg, col_reg}<16'b1000001101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000001101100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001101100100) && ({row_reg, col_reg}<16'b1000001101100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001101100111) && ({row_reg, col_reg}<16'b1000001101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001101101010) && ({row_reg, col_reg}<16'b1000001101101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001101101101) && ({row_reg, col_reg}<16'b1000001101110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000001101110111) && ({row_reg, col_reg}<16'b1000001101111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001101111100) && ({row_reg, col_reg}<16'b1000001101111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000001101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001110000000) && ({row_reg, col_reg}<16'b1000001110000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001110000101) && ({row_reg, col_reg}<16'b1000001110000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001110000111) && ({row_reg, col_reg}<16'b1000001110010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000001110010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001110010100) && ({row_reg, col_reg}<16'b1000001110011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001110011000) && ({row_reg, col_reg}<16'b1000001110011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001110011011) && ({row_reg, col_reg}<16'b1000001110011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001110011101) && ({row_reg, col_reg}<16'b1000001110100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001110100000) && ({row_reg, col_reg}<16'b1000001110100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001110100010) && ({row_reg, col_reg}<16'b1000001110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000001110101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000001110101100) && ({row_reg, col_reg}<16'b1000001110101110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000001110101110) && ({row_reg, col_reg}<16'b1000001110110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000001110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000001110110110) && ({row_reg, col_reg}<16'b1000001110111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000001110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001110111011) && ({row_reg, col_reg}<16'b1000001110111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000001110111110) && ({row_reg, col_reg}<16'b1000001111000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001111000010) && ({row_reg, col_reg}<16'b1000001111000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000001111000110) && ({row_reg, col_reg}<16'b1000001111001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000001111001010) && ({row_reg, col_reg}<16'b1000001111001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000001111001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001111001101) && ({row_reg, col_reg}<16'b1000001111010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000001111010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000001111010100) && ({row_reg, col_reg}<16'b1000001111010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000001111010111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000001111011000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000001111011001) && ({row_reg, col_reg}<16'b1000001111011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000001111011011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000001111011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000001111011101) && ({row_reg, col_reg}<16'b1000001111100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000001111100110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000001111100111) && ({row_reg, col_reg}<16'b1000001111101110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001111101110) && ({row_reg, col_reg}<16'b1000001111110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001111110001) && ({row_reg, col_reg}<16'b1000001111110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000001111110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001111110100) && ({row_reg, col_reg}<16'b1000001111110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000001111110110) && ({row_reg, col_reg}<16'b1000001111111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000001111111000) && ({row_reg, col_reg}<16'b1000001111111101)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}>=16'b1000001111111101) && ({row_reg, col_reg}<16'b1000010000000000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000010000000000) && ({row_reg, col_reg}<16'b1000010000000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010000000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000010000000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010000000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000010000000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000010000000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010000001000) && ({row_reg, col_reg}<16'b1000010000001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000010000001010) && ({row_reg, col_reg}<16'b1000010000001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000010000001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010000001101) && ({row_reg, col_reg}<16'b1000010000001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000010000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010000010000) && ({row_reg, col_reg}<16'b1000010000010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000010000010100) && ({row_reg, col_reg}<16'b1000010001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000010001100011) && ({row_reg, col_reg}<16'b1000010001101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010001101010) && ({row_reg, col_reg}<16'b1000010001101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010001101101) && ({row_reg, col_reg}<16'b1000010001110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010001110100) && ({row_reg, col_reg}<16'b1000010001110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000010001110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000010001110111) && ({row_reg, col_reg}<16'b1000010001111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010001111100) && ({row_reg, col_reg}<16'b1000010001111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000010001111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000010001111111) && ({row_reg, col_reg}<16'b1000010010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010010000001) && ({row_reg, col_reg}<16'b1000010010010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010010010010) && ({row_reg, col_reg}<16'b1000010010010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010010010101) && ({row_reg, col_reg}<16'b1000010010011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010010011000) && ({row_reg, col_reg}<16'b1000010010011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010010011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010010011101) && ({row_reg, col_reg}<16'b1000010010100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010010100011) && ({row_reg, col_reg}<16'b1000010010100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010010100101) && ({row_reg, col_reg}<16'b1000010010101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010010101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000010010101010) && ({row_reg, col_reg}<16'b1000010010101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010010101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000010010101101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000010010101110) && ({row_reg, col_reg}<16'b1000010010110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000010010110011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000010010110100) && ({row_reg, col_reg}<16'b1000010010110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000010010110111) && ({row_reg, col_reg}<16'b1000010010111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000010010111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010010111011) && ({row_reg, col_reg}<16'b1000010010111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000010010111101) && ({row_reg, col_reg}<16'b1000010011000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000010011000010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000010011000011) && ({row_reg, col_reg}<16'b1000010011000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000010011000111) && ({row_reg, col_reg}<16'b1000010011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010011001010) && ({row_reg, col_reg}<16'b1000010011001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000010011001110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000010011001111) && ({row_reg, col_reg}<16'b1000010011010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010011010001) && ({row_reg, col_reg}<16'b1000010011010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010011010111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010011011000) && ({row_reg, col_reg}<16'b1000010011011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000010011011110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000010011011111) && ({row_reg, col_reg}<16'b1000010011100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000010011100101) && ({row_reg, col_reg}<16'b1000010011100111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000010011100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000010011101000) && ({row_reg, col_reg}<16'b1000010011101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010011101010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000010011101011) && ({row_reg, col_reg}<16'b1000010011110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000010011110001) && ({row_reg, col_reg}<16'b1000010011110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010011110011) && ({row_reg, col_reg}<16'b1000010011110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010011110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000010011111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010011111001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000010011111010) && ({row_reg, col_reg}<16'b1000010011111110)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}>=16'b1000010011111110) && ({row_reg, col_reg}<16'b1000010100000000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000010100000000) && ({row_reg, col_reg}<16'b1000010100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010100000010) && ({row_reg, col_reg}<16'b1000010100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010100000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010100000111) && ({row_reg, col_reg}<16'b1000010100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000010100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010100001010) && ({row_reg, col_reg}<16'b1000010100001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010100001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010100001111) && ({row_reg, col_reg}<16'b1000010100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010100010001) && ({row_reg, col_reg}<16'b1000010100010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000010100010100) && ({row_reg, col_reg}<16'b1000010101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000010101100011) && ({row_reg, col_reg}<16'b1000010101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010101101010) && ({row_reg, col_reg}<16'b1000010101101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010101101101) && ({row_reg, col_reg}<16'b1000010101110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010101110101) && ({row_reg, col_reg}<16'b1000010101110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010101110111) && ({row_reg, col_reg}<16'b1000010101111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010101111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000010101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010101111100) && ({row_reg, col_reg}<16'b1000010101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000010101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000010101111111) && ({row_reg, col_reg}<16'b1000010110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010110000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010110000010) && ({row_reg, col_reg}<16'b1000010110001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010110001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010110001010) && ({row_reg, col_reg}<16'b1000010110001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010110001101) && ({row_reg, col_reg}<16'b1000010110010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010110010000) && ({row_reg, col_reg}<16'b1000010110011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010110011000) && ({row_reg, col_reg}<16'b1000010110011011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000010110011011) && ({row_reg, col_reg}<16'b1000010110100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010110100010) && ({row_reg, col_reg}<16'b1000010110100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010110100110) && ({row_reg, col_reg}<16'b1000010110101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000010110101000) && ({row_reg, col_reg}<16'b1000010110101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000010110101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010110101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000010110101110) && ({row_reg, col_reg}<16'b1000010110110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000010110110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000010110110001) && ({row_reg, col_reg}<16'b1000010110110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010110110011) && ({row_reg, col_reg}<16'b1000010110111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000010110111010) && ({row_reg, col_reg}<16'b1000010110111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000010110111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000010110111101) && ({row_reg, col_reg}<16'b1000010111000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010111000010) && ({row_reg, col_reg}<16'b1000010111000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000010111000101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000010111000110) && ({row_reg, col_reg}<16'b1000010111001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000010111001011) && ({row_reg, col_reg}<16'b1000010111001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000010111001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000010111010000) && ({row_reg, col_reg}<16'b1000010111010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010111010010) && ({row_reg, col_reg}<16'b1000010111010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010111010100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010111010101) && ({row_reg, col_reg}<16'b1000010111011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000010111011010) && ({row_reg, col_reg}<16'b1000010111011100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010111011100) && ({row_reg, col_reg}<16'b1000010111011111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000010111011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010111100000) && ({row_reg, col_reg}<16'b1000010111100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000010111100010) && ({row_reg, col_reg}<16'b1000010111101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000010111101000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010111101001) && ({row_reg, col_reg}<16'b1000010111101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000010111101101) && ({row_reg, col_reg}<16'b1000010111110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010111110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000010111110011) && ({row_reg, col_reg}<16'b1000010111111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000010111111000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010111111001) && ({row_reg, col_reg}<16'b1000010111111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000010111111011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000010111111100) && ({row_reg, col_reg}<16'b1000010111111110)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}>=16'b1000010111111110) && ({row_reg, col_reg}<16'b1000011000000000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000011000000000) && ({row_reg, col_reg}<16'b1000011000000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011000000010) && ({row_reg, col_reg}<16'b1000011000000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011000000111) && ({row_reg, col_reg}<16'b1000011000001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011000001011) && ({row_reg, col_reg}<16'b1000011000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011000001111) && ({row_reg, col_reg}<16'b1000011000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011000010001) && ({row_reg, col_reg}<16'b1000011000010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000011000010100) && ({row_reg, col_reg}<16'b1000011001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000011001100011) && ({row_reg, col_reg}<16'b1000011001100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011001100101) && ({row_reg, col_reg}<16'b1000011001101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011001101001) && ({row_reg, col_reg}<16'b1000011001101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011001101101) && ({row_reg, col_reg}<16'b1000011001110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011001110110) && ({row_reg, col_reg}<16'b1000011001111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011001111000) && ({row_reg, col_reg}<16'b1000011001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000011001111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000011001111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000011001111101) && ({row_reg, col_reg}<16'b1000011001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000011001111111) && ({row_reg, col_reg}<16'b1000011010000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000011010000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011010000010) && ({row_reg, col_reg}<16'b1000011010001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000011010001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011010001010) && ({row_reg, col_reg}<16'b1000011010001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011010001101) && ({row_reg, col_reg}<16'b1000011010001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011010001111) && ({row_reg, col_reg}<16'b1000011010011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011010011001) && ({row_reg, col_reg}<16'b1000011010011011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011010011011) && ({row_reg, col_reg}<16'b1000011010100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011010100001) && ({row_reg, col_reg}<16'b1000011010100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000011010100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000011010100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011010100111) && ({row_reg, col_reg}<16'b1000011010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011010101010) && ({row_reg, col_reg}<16'b1000011010101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000011010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000011010101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000011010101111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000011010110000) && ({row_reg, col_reg}<16'b1000011010110010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000011010110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000011010110011) && ({row_reg, col_reg}<16'b1000011010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011010110101) && ({row_reg, col_reg}<16'b1000011010111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000011010111100) && ({row_reg, col_reg}<16'b1000011010111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000011010111111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1000011011000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000011011000001) && ({row_reg, col_reg}<16'b1000011011000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011011000101) && ({row_reg, col_reg}<16'b1000011011001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000011011001000) && ({row_reg, col_reg}<16'b1000011011001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011011001011) && ({row_reg, col_reg}<16'b1000011011010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000011011010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011011010001) && ({row_reg, col_reg}<16'b1000011011010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000011011010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000011011010100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000011011010101) && ({row_reg, col_reg}<16'b1000011011011001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000011011011001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000011011011010) && ({row_reg, col_reg}<16'b1000011011011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000011011011100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000011011011101) && ({row_reg, col_reg}<16'b1000011011100000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000011011100000) && ({row_reg, col_reg}<16'b1000011011100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000011011100010) && ({row_reg, col_reg}<16'b1000011011101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000011011101101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000011011101110) && ({row_reg, col_reg}<16'b1000011011110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000011011110101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000011011110110) && ({row_reg, col_reg}<16'b1000011011111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000011011111011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000011011111100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000011011111101)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}>=16'b1000011011111110) && ({row_reg, col_reg}<16'b1000011100000000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000011100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011100000001) && ({row_reg, col_reg}<16'b1000011100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000011100000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000011100000111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000011100001000) && ({row_reg, col_reg}<16'b1000011100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011100001100) && ({row_reg, col_reg}<16'b1000011100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011100001111) && ({row_reg, col_reg}<16'b1000011100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011100010001) && ({row_reg, col_reg}<16'b1000011100010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000011100010100) && ({row_reg, col_reg}<16'b1000011101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000011101100011) && ({row_reg, col_reg}<16'b1000011101100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011101100101) && ({row_reg, col_reg}<16'b1000011101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011101101010) && ({row_reg, col_reg}<16'b1000011101101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011101101101) && ({row_reg, col_reg}<16'b1000011101110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011101110110) && ({row_reg, col_reg}<16'b1000011101111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011101111000) && ({row_reg, col_reg}<16'b1000011101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011101111011) && ({row_reg, col_reg}<16'b1000011101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000011101111111) && ({row_reg, col_reg}<16'b1000011110001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011110001000) && ({row_reg, col_reg}<16'b1000011110001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000011110001010) && ({row_reg, col_reg}<16'b1000011110001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011110001100) && ({row_reg, col_reg}<16'b1000011110001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000011110001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011110001111) && ({row_reg, col_reg}<16'b1000011110010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011110010010) && ({row_reg, col_reg}<16'b1000011110100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000011110100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011110100110) && ({row_reg, col_reg}<16'b1000011110101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011110101010) && ({row_reg, col_reg}<16'b1000011110101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000011110101101) && ({row_reg, col_reg}<16'b1000011110110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011110110000) && ({row_reg, col_reg}<16'b1000011110110011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000011110110011) && ({row_reg, col_reg}<16'b1000011110110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000011110110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000011110110111) && ({row_reg, col_reg}<16'b1000011110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000011110111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011110111011) && ({row_reg, col_reg}<16'b1000011110111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000011110111111) && ({row_reg, col_reg}<16'b1000011111000001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000011111000001) && ({row_reg, col_reg}<16'b1000011111000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000011111000011) && ({row_reg, col_reg}<16'b1000011111000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000011111000111) && ({row_reg, col_reg}<16'b1000011111001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000011111001001) && ({row_reg, col_reg}<16'b1000011111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000011111010001) && ({row_reg, col_reg}<16'b1000011111010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000011111010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000011111010100) && ({row_reg, col_reg}<16'b1000011111011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000011111011000) && ({row_reg, col_reg}<16'b1000011111011010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000011111011010) && ({row_reg, col_reg}<16'b1000011111011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000011111011101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000011111011110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000011111011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000011111100000) && ({row_reg, col_reg}<16'b1000011111100010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000011111100010) && ({row_reg, col_reg}<16'b1000011111100101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000011111100101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000011111100110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000011111100111) && ({row_reg, col_reg}<16'b1000011111101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000011111101001) && ({row_reg, col_reg}<16'b1000011111101100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000011111101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000011111101101) && ({row_reg, col_reg}<16'b1000011111110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000011111110011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000011111110100) && ({row_reg, col_reg}<16'b1000011111111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000011111111010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000011111111011) && ({row_reg, col_reg}<16'b1000011111111101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000011111111101) && ({row_reg, col_reg}<16'b1000011111111111)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}==16'b1000011111111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000100000000000) && ({row_reg, col_reg}<16'b1000100000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100000000110) && ({row_reg, col_reg}<16'b1000100000001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000100000001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000100000001001) && ({row_reg, col_reg}<16'b1000100000001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100000001101) && ({row_reg, col_reg}<16'b1000100000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100000010001) && ({row_reg, col_reg}<16'b1000100000010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100000010100) && ({row_reg, col_reg}<16'b1000100001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000100001100011) && ({row_reg, col_reg}<16'b1000100001100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100001100110) && ({row_reg, col_reg}<16'b1000100001101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100001101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100001101100) && ({row_reg, col_reg}<16'b1000100001110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100001110111) && ({row_reg, col_reg}<16'b1000100001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100001111011) && ({row_reg, col_reg}<16'b1000100001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100001111111) && ({row_reg, col_reg}<16'b1000100010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100010000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100010000011) && ({row_reg, col_reg}<16'b1000100010000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100010000111) && ({row_reg, col_reg}<16'b1000100010001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100010001001) && ({row_reg, col_reg}<16'b1000100010001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100010001011) && ({row_reg, col_reg}<16'b1000100010001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100010001101) && ({row_reg, col_reg}<16'b1000100010010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100010010011) && ({row_reg, col_reg}<16'b1000100010011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100010011100) && ({row_reg, col_reg}<16'b1000100010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100010011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100010100000) && ({row_reg, col_reg}<16'b1000100010101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100010101000) && ({row_reg, col_reg}<16'b1000100010101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100010101010) && ({row_reg, col_reg}<16'b1000100010101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100010101100) && ({row_reg, col_reg}<16'b1000100010101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100010101110) && ({row_reg, col_reg}<16'b1000100010110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100010110011) && ({row_reg, col_reg}<16'b1000100010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000100010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000100010110110) && ({row_reg, col_reg}<16'b1000100011000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000100011000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000100011000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000100011000011) && ({row_reg, col_reg}<16'b1000100011000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000100011000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000100011000111) && ({row_reg, col_reg}<16'b1000100011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100011001010) && ({row_reg, col_reg}<16'b1000100011010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000100011010101) && ({row_reg, col_reg}<16'b1000100011010111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1000100011010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000100011011000) && ({row_reg, col_reg}<16'b1000100011011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000100011011011) && ({row_reg, col_reg}<16'b1000100011011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000100011011101) && ({row_reg, col_reg}<16'b1000100011100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100011100001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000100011100010) && ({row_reg, col_reg}<16'b1000100011100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100011100110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000100011100111) && ({row_reg, col_reg}<16'b1000100011101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000100011101001) && ({row_reg, col_reg}<16'b1000100011101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100011101100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000100011101101) && ({row_reg, col_reg}<16'b1000100011110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000100011110010) && ({row_reg, col_reg}<16'b1000100011111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000100011111010) && ({row_reg, col_reg}<16'b1000100011111100)) color_data = 12'b010000100001;

		if(({row_reg, col_reg}>=16'b1000100011111100) && ({row_reg, col_reg}<16'b1000100100000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000100100000000) && ({row_reg, col_reg}<16'b1000100100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100100000110) && ({row_reg, col_reg}<16'b1000100100001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000100100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000100100001010) && ({row_reg, col_reg}<16'b1000100100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000100100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100100001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000100100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100100010000) && ({row_reg, col_reg}<16'b1000100100010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100100010100) && ({row_reg, col_reg}<16'b1000100101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000100101100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100101100100) && ({row_reg, col_reg}<16'b1000100101100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100101100110) && ({row_reg, col_reg}<16'b1000100101110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100101110111) && ({row_reg, col_reg}<16'b1000100101111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000100101111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100101111011) && ({row_reg, col_reg}<16'b1000100101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100101111111) && ({row_reg, col_reg}<16'b1000100110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100110000001) && ({row_reg, col_reg}<16'b1000100110000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100110000011) && ({row_reg, col_reg}<16'b1000100110000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100110000111) && ({row_reg, col_reg}<16'b1000100110001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100110001001) && ({row_reg, col_reg}<16'b1000100110001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100110001111) && ({row_reg, col_reg}<16'b1000100110011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100110011011) && ({row_reg, col_reg}<16'b1000100110011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100110011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000100110011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100110011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100110100000) && ({row_reg, col_reg}<16'b1000100110100011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100110100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100110100100) && ({row_reg, col_reg}<16'b1000100110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000100110101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100110101010) && ({row_reg, col_reg}<16'b1000100110101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100110101100) && ({row_reg, col_reg}<16'b1000100110101111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000100110101111) && ({row_reg, col_reg}<16'b1000100110110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000100110110011) && ({row_reg, col_reg}<16'b1000100110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000100110110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000100110110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000100110110111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000100110111000) && ({row_reg, col_reg}<16'b1000100111000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000100111000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000100111000010) && ({row_reg, col_reg}<16'b1000100111000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000100111000100) && ({row_reg, col_reg}<16'b1000100111000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000100111000110) && ({row_reg, col_reg}<16'b1000100111001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000100111001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000100111001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000100111001011) && ({row_reg, col_reg}<16'b1000100111001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000100111001111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1000100111010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000100111010001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000100111010010) && ({row_reg, col_reg}<16'b1000100111010111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000100111010111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000100111011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000100111011001) && ({row_reg, col_reg}<16'b1000100111011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100111011011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000100111011100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000100111011101) && ({row_reg, col_reg}<16'b1000100111100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000100111100001) && ({row_reg, col_reg}<16'b1000100111100011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000100111100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100111100100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000100111100101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000100111100110) && ({row_reg, col_reg}<16'b1000100111101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000100111101001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000100111101010) && ({row_reg, col_reg}<16'b1000100111101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100111101100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000100111101101) && ({row_reg, col_reg}<16'b1000100111110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000100111110010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000100111110011) && ({row_reg, col_reg}<16'b1000100111111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000100111111011)) color_data = 12'b010000110001;

		if(({row_reg, col_reg}>=16'b1000100111111100) && ({row_reg, col_reg}<16'b1000101000000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000101000000000) && ({row_reg, col_reg}<16'b1000101000000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000101000000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101000000100) && ({row_reg, col_reg}<16'b1000101000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101000000110) && ({row_reg, col_reg}<16'b1000101000001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000101000001010) && ({row_reg, col_reg}<16'b1000101000001100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000101000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000101000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000101000001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000101000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101000010000) && ({row_reg, col_reg}<16'b1000101000010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101000010100) && ({row_reg, col_reg}<16'b1000101001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000101001100011) && ({row_reg, col_reg}<16'b1000101001100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101001100101) && ({row_reg, col_reg}<16'b1000101001111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000101001111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000101001111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101001111011) && ({row_reg, col_reg}<16'b1000101001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101001111111) && ({row_reg, col_reg}<16'b1000101010001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101010001110) && ({row_reg, col_reg}<16'b1000101010011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101010011100) && ({row_reg, col_reg}<16'b1000101010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101010011111) && ({row_reg, col_reg}<16'b1000101010100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101010100001) && ({row_reg, col_reg}<16'b1000101010100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000101010100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101010100110) && ({row_reg, col_reg}<16'b1000101010110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101010110000) && ({row_reg, col_reg}<16'b1000101010110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000101010110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101010110011) && ({row_reg, col_reg}<16'b1000101010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000101010110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000101010110111) && ({row_reg, col_reg}<16'b1000101010111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101010111001) && ({row_reg, col_reg}<16'b1000101010111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000101010111011) && ({row_reg, col_reg}<16'b1000101010111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101010111110) && ({row_reg, col_reg}<16'b1000101011000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000101011000001) && ({row_reg, col_reg}<16'b1000101011000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101011000011) && ({row_reg, col_reg}<16'b1000101011000111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000101011000111) && ({row_reg, col_reg}<16'b1000101011001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000101011001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000101011001010) && ({row_reg, col_reg}<16'b1000101011001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101011001100) && ({row_reg, col_reg}<16'b1000101011001111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000101011001111) && ({row_reg, col_reg}<16'b1000101011010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101011010011) && ({row_reg, col_reg}<16'b1000101011010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000101011010101) && ({row_reg, col_reg}<16'b1000101011011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101011011000) && ({row_reg, col_reg}<16'b1000101011011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000101011011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101011011011) && ({row_reg, col_reg}<16'b1000101011100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000101011100001) && ({row_reg, col_reg}<16'b1000101011100101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000101011100101) && ({row_reg, col_reg}<16'b1000101011101001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000101011101001) && ({row_reg, col_reg}<16'b1000101011101011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000101011101011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000101011101100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000101011101101) && ({row_reg, col_reg}<16'b1000101011110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000101011110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000101011110011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000101011110100) && ({row_reg, col_reg}<16'b1000101011110110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000101011110110) && ({row_reg, col_reg}<16'b1000101011111000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000101011111000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000101011111001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000101011111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000101011111011)) color_data = 12'b010000110001;

		if(({row_reg, col_reg}>=16'b1000101011111100) && ({row_reg, col_reg}<16'b1000101100000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000101100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101100000001) && ({row_reg, col_reg}<16'b1000101100000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000101100000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101100000100) && ({row_reg, col_reg}<16'b1000101100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101100000110) && ({row_reg, col_reg}<16'b1000101100001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000101100001011) && ({row_reg, col_reg}<16'b1000101100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101100001101) && ({row_reg, col_reg}<16'b1000101100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101100010001) && ({row_reg, col_reg}<16'b1000101100010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101100010100) && ({row_reg, col_reg}<16'b1000101101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000101101100011) && ({row_reg, col_reg}<16'b1000101101100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101101100101) && ({row_reg, col_reg}<16'b1000101101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101101101010) && ({row_reg, col_reg}<16'b1000101101110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101101110000) && ({row_reg, col_reg}<16'b1000101101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101101111011) && ({row_reg, col_reg}<16'b1000101101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101101111111) && ({row_reg, col_reg}<16'b1000101110001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101110001101) && ({row_reg, col_reg}<16'b1000101110011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101110011101) && ({row_reg, col_reg}<16'b1000101110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101110011111) && ({row_reg, col_reg}<16'b1000101110100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000101110100010) && ({row_reg, col_reg}<16'b1000101110110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000101110110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000101110110010) && ({row_reg, col_reg}<16'b1000101110110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000101110110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000101110110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101110111000) && ({row_reg, col_reg}<16'b1000101110111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000101110111010) && ({row_reg, col_reg}<16'b1000101110111110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101110111110) && ({row_reg, col_reg}<16'b1000101111000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000101111000001) && ({row_reg, col_reg}<16'b1000101111000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000101111000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000101111000100) && ({row_reg, col_reg}<16'b1000101111000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101111000111) && ({row_reg, col_reg}<16'b1000101111001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000101111001010) && ({row_reg, col_reg}<16'b1000101111001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000101111001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000101111001101) && ({row_reg, col_reg}<16'b1000101111010000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000101111010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000101111010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000101111010010) && ({row_reg, col_reg}<16'b1000101111010100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101111010100) && ({row_reg, col_reg}<16'b1000101111010111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000101111010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000101111011000) && ({row_reg, col_reg}<16'b1000101111011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000101111011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000101111011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000101111011100) && ({row_reg, col_reg}<16'b1000101111011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000101111011111) && ({row_reg, col_reg}<16'b1000101111100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000101111100010) && ({row_reg, col_reg}<16'b1000101111100101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000101111100101) && ({row_reg, col_reg}<16'b1000101111101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000101111101000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000101111101001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000101111101010) && ({row_reg, col_reg}<16'b1000101111101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000101111101100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000101111101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000101111101110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000101111101111) && ({row_reg, col_reg}<16'b1000101111110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000101111110010) && ({row_reg, col_reg}<16'b1000101111110110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000101111110110) && ({row_reg, col_reg}<16'b1000101111111010)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}>=16'b1000101111111010) && ({row_reg, col_reg}<16'b1000110000000000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110000000000) && ({row_reg, col_reg}<16'b1000110000000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110000000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000110000000100) && ({row_reg, col_reg}<16'b1000110000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110000000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110000000111) && ({row_reg, col_reg}<16'b1000110000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000110000001001) && ({row_reg, col_reg}<16'b1000110000001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000110000001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000110000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110000001110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000110000001111) && ({row_reg, col_reg}<16'b1000110000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110000010001) && ({row_reg, col_reg}<16'b1000110000010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000110000010011) && ({row_reg, col_reg}<16'b1000110001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000110001100011) && ({row_reg, col_reg}<16'b1000110001101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110001101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000110001101011)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==16'b1000110001101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000110001101101) && ({row_reg, col_reg}<16'b1000110001110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110001110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000110001111000) && ({row_reg, col_reg}<16'b1000110001111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110001111011) && ({row_reg, col_reg}<16'b1000110001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000110001111111) && ({row_reg, col_reg}<16'b1000110010000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110010000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000110010001000) && ({row_reg, col_reg}<16'b1000110010001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110010001100) && ({row_reg, col_reg}<16'b1000110010010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110010010010) && ({row_reg, col_reg}<16'b1000110010010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110010010101) && ({row_reg, col_reg}<16'b1000110010011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110010011000) && ({row_reg, col_reg}<16'b1000110010011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110010011100) && ({row_reg, col_reg}<16'b1000110010011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000110010011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110010011111) && ({row_reg, col_reg}<16'b1000110010100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110010100011) && ({row_reg, col_reg}<16'b1000110010110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110010110011) && ({row_reg, col_reg}<16'b1000110010110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000110010110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000110010110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000110010111000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110010111001) && ({row_reg, col_reg}<16'b1000110010111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1000110010111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110011000000) && ({row_reg, col_reg}<16'b1000110011000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000110011000011) && ({row_reg, col_reg}<16'b1000110011000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110011000101) && ({row_reg, col_reg}<16'b1000110011000111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000110011000111) && ({row_reg, col_reg}<16'b1000110011001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110011001100) && ({row_reg, col_reg}<16'b1000110011001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000110011001110) && ({row_reg, col_reg}<16'b1000110011010000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000110011010000) && ({row_reg, col_reg}<16'b1000110011010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110011010101) && ({row_reg, col_reg}<16'b1000110011010111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000110011010111) && ({row_reg, col_reg}<16'b1000110011011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110011011010) && ({row_reg, col_reg}<16'b1000110011011111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000110011011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110011100000) && ({row_reg, col_reg}<16'b1000110011100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000110011100101) && ({row_reg, col_reg}<16'b1000110011101000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000110011101000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000110011101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000110011101010) && ({row_reg, col_reg}<16'b1000110011101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000110011101111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110011110000) && ({row_reg, col_reg}<16'b1000110011110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110011110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110011110011) && ({row_reg, col_reg}<16'b1000110011110101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000110011110101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110011110110) && ({row_reg, col_reg}<16'b1000110011111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110011111000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000110011111001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000110011111010) && ({row_reg, col_reg}<16'b1000110011111111)) color_data = 12'b010000100001;

		if(({row_reg, col_reg}==16'b1000110011111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000110100000000) && ({row_reg, col_reg}<16'b1000110100000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110100000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000110100000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110100000101) && ({row_reg, col_reg}<16'b1000110100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110100001001) && ({row_reg, col_reg}<16'b1000110100001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000110100001011) && ({row_reg, col_reg}<16'b1000110100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110100001101) && ({row_reg, col_reg}<16'b1000110100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000110100001111) && ({row_reg, col_reg}<16'b1000110100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110100010001) && ({row_reg, col_reg}<16'b1000110100010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000110100010011) && ({row_reg, col_reg}<16'b1000110101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000110101100011) && ({row_reg, col_reg}<16'b1000110101101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110101101001) && ({row_reg, col_reg}<16'b1000110101101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000110101101011) && ({row_reg, col_reg}<16'b1000110101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000110101101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000110101101110) && ({row_reg, col_reg}<16'b1000110101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110101111011) && ({row_reg, col_reg}<16'b1000110101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000110101111111) && ({row_reg, col_reg}<16'b1000110110000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110110000011) && ({row_reg, col_reg}<16'b1000110110000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110110000101) && ({row_reg, col_reg}<16'b1000110110001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110110001010) && ({row_reg, col_reg}<16'b1000110110010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110110010010) && ({row_reg, col_reg}<16'b1000110110010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110110010101) && ({row_reg, col_reg}<16'b1000110110011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110110011000) && ({row_reg, col_reg}<16'b1000110110011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000110110011100) && ({row_reg, col_reg}<16'b1000110110101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000110110101111) && ({row_reg, col_reg}<16'b1000110110111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110110111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000110110111001) && ({row_reg, col_reg}<16'b1000110111000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000110111000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000110111000001) && ({row_reg, col_reg}<16'b1000110111001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000110111001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000110111001010) && ({row_reg, col_reg}<16'b1000110111001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110111001110) && ({row_reg, col_reg}<16'b1000110111010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1000110111010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000110111010011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000110111010100) && ({row_reg, col_reg}<16'b1000110111010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000110111010110) && ({row_reg, col_reg}<16'b1000110111011101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000110111011101) && ({row_reg, col_reg}<16'b1000110111011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000110111011111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000110111100000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000110111100001) && ({row_reg, col_reg}<16'b1000110111100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110111100101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000110111100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000110111100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000110111101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110111101001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110111101010) && ({row_reg, col_reg}<16'b1000110111101111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000110111101111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110111110000) && ({row_reg, col_reg}<16'b1000110111110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000110111110011) && ({row_reg, col_reg}<16'b1000110111110101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000110111110101) && ({row_reg, col_reg}<16'b1000110111110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110111110111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110111111000) && ({row_reg, col_reg}<16'b1000110111111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000110111111010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000110111111011) && ({row_reg, col_reg}<16'b1000110111111110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000110111111110)) color_data = 12'b010000110001;

		if(({row_reg, col_reg}==16'b1000110111111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=16'b1000111000000000) && ({row_reg, col_reg}<16'b1000111000000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000111000000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000111000000100) && ({row_reg, col_reg}<16'b1000111000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000111000000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000111000000111) && ({row_reg, col_reg}<16'b1000111000001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000111000001001) && ({row_reg, col_reg}<16'b1000111000001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000111000001011) && ({row_reg, col_reg}<16'b1000111000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111000001101) && ({row_reg, col_reg}<16'b1000111000001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000111000001111) && ({row_reg, col_reg}<16'b1000111000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111000010001) && ({row_reg, col_reg}<16'b1000111000010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000111000010100) && ({row_reg, col_reg}<16'b1000111001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000111001100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111001100100) && ({row_reg, col_reg}<16'b1000111001101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111001101000) && ({row_reg, col_reg}<16'b1000111001101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000111001101010) && ({row_reg, col_reg}<16'b1000111001101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000111001101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000111001101110) && ({row_reg, col_reg}<16'b1000111001111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111001111010) && ({row_reg, col_reg}<16'b1000111001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000111001111111) && ({row_reg, col_reg}<16'b1000111010000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111010000011) && ({row_reg, col_reg}<16'b1000111010000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111010000110) && ({row_reg, col_reg}<16'b1000111010001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111010001001) && ({row_reg, col_reg}<16'b1000111010010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000111010010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111010010100) && ({row_reg, col_reg}<16'b1000111010010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111010010110) && ({row_reg, col_reg}<16'b1000111010011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000111010011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000111010011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111010011011) && ({row_reg, col_reg}<16'b1000111010101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111010101111) && ({row_reg, col_reg}<16'b1000111010111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000111010111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000111010111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000111010111011) && ({row_reg, col_reg}<16'b1000111011000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000111011000001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000111011000010) && ({row_reg, col_reg}<16'b1000111011001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000111011001110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000111011001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000111011010000)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==16'b1000111011010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1000111011010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000111011010011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1000111011010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000111011010101) && ({row_reg, col_reg}<16'b1000111011010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111011010111) && ({row_reg, col_reg}<16'b1000111011011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000111011011010) && ({row_reg, col_reg}<16'b1000111011011101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000111011011101) && ({row_reg, col_reg}<16'b1000111011100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000111011100000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000111011100001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000111011100010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111011100011) && ({row_reg, col_reg}<16'b1000111011100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111011100101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000111011100110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000111011100111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==16'b1000111011101000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000111011101001) && ({row_reg, col_reg}<16'b1000111011101110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000111011101110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000111011101111) && ({row_reg, col_reg}<16'b1000111011110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1000111011110011) && ({row_reg, col_reg}<16'b1000111011110101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000111011110101) && ({row_reg, col_reg}<16'b1000111011111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111011111000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000111011111001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000111011111010) && ({row_reg, col_reg}<16'b1000111011111110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111011111110)) color_data = 12'b010000100001;

		if(({row_reg, col_reg}==16'b1000111011111111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1000111100000000) && ({row_reg, col_reg}<16'b1000111100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111100000110) && ({row_reg, col_reg}<16'b1000111100001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000111100001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000111100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000111100001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111100001101) && ({row_reg, col_reg}<16'b1000111100001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000111100001111) && ({row_reg, col_reg}<16'b1000111100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111100010001) && ({row_reg, col_reg}<16'b1000111100010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000111100010100) && ({row_reg, col_reg}<16'b1000111101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000111101100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1000111101100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111101100101) && ({row_reg, col_reg}<16'b1000111101101000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000111101101000) && ({row_reg, col_reg}<16'b1000111101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1000111101101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000111101101110) && ({row_reg, col_reg}<16'b1000111101111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111101111010) && ({row_reg, col_reg}<16'b1000111101111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000111101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1000111110000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1000111110000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111110000010) && ({row_reg, col_reg}<16'b1000111110000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111110000110) && ({row_reg, col_reg}<16'b1000111110001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111110001001) && ({row_reg, col_reg}<16'b1000111110001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111110001011) && ({row_reg, col_reg}<16'b1000111110010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111110010011) && ({row_reg, col_reg}<16'b1000111110010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111110010101) && ({row_reg, col_reg}<16'b1000111110011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111110011000) && ({row_reg, col_reg}<16'b1000111110101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1000111110101111) && ({row_reg, col_reg}<16'b1000111110110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111110110111) && ({row_reg, col_reg}<16'b1000111110111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1000111110111001) && ({row_reg, col_reg}<16'b1000111110111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111110111011) && ({row_reg, col_reg}<16'b1000111110111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000111110111101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000111110111110) && ({row_reg, col_reg}<16'b1000111111000001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000111111000001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1000111111000010) && ({row_reg, col_reg}<16'b1000111111000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111111000100) && ({row_reg, col_reg}<16'b1000111111000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000111111000111) && ({row_reg, col_reg}<16'b1000111111001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111111001010) && ({row_reg, col_reg}<16'b1000111111001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1000111111001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111111001101) && ({row_reg, col_reg}<16'b1000111111001111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1000111111001111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000111111010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1000111111010001) && ({row_reg, col_reg}<16'b1000111111011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1000111111011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1000111111011100) && ({row_reg, col_reg}<16'b1000111111011111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1000111111011111) && ({row_reg, col_reg}<16'b1000111111100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1000111111100010) && ({row_reg, col_reg}<16'b1000111111100100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1000111111100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1000111111100101) && ({row_reg, col_reg}<16'b1000111111101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111111101000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000111111101001) && ({row_reg, col_reg}<16'b1000111111101101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1000111111101101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==16'b1000111111101110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1000111111101111) && ({row_reg, col_reg}<16'b1000111111110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1000111111110100)) color_data = 12'b010000100001;

		if(({row_reg, col_reg}>=16'b1000111111110101) && ({row_reg, col_reg}<16'b1001000000000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001000000000000) && ({row_reg, col_reg}<16'b1001000000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000000000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001000000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000000000111) && ({row_reg, col_reg}<16'b1001000000001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001000000001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000000001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000000001100) && ({row_reg, col_reg}<16'b1001000000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000000010001) && ({row_reg, col_reg}<16'b1001000000010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001000000010100) && ({row_reg, col_reg}<16'b1001000001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001000001100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001000001100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000001100101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001000001100110) && ({row_reg, col_reg}<16'b1001000001101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001000001101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001000001101101) && ({row_reg, col_reg}<16'b1001000001111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000001111010) && ({row_reg, col_reg}<16'b1001000001111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001000001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000010000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001000010000001) && ({row_reg, col_reg}<16'b1001000010000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000010000011) && ({row_reg, col_reg}<16'b1001000010000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001000010000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000010001000) && ({row_reg, col_reg}<16'b1001000010001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000010001011) && ({row_reg, col_reg}<16'b1001000010010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000010010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001000010010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000010010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000010010100) && ({row_reg, col_reg}<16'b1001000010010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000010010111) && ({row_reg, col_reg}<16'b1001000010100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000010100010) && ({row_reg, col_reg}<16'b1001000010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000010100100) && ({row_reg, col_reg}<16'b1001000010101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000010101111) && ({row_reg, col_reg}<16'b1001000010110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000010110011) && ({row_reg, col_reg}<16'b1001000010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001000010110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000010110110) && ({row_reg, col_reg}<16'b1001000010111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001000010111001) && ({row_reg, col_reg}<16'b1001000010111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000010111011) && ({row_reg, col_reg}<16'b1001000010111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001000010111101) && ({row_reg, col_reg}<16'b1001000011000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001000011000001) && ({row_reg, col_reg}<16'b1001000011000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000011000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001000011000101) && ({row_reg, col_reg}<16'b1001000011001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000011001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001000011001010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=16'b1001000011001011) && ({row_reg, col_reg}<16'b1001000011001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001000011001101)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}>=16'b1001000011001110) && ({row_reg, col_reg}<16'b1001000011010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001000011010000) && ({row_reg, col_reg}<16'b1001000011010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000011010010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001000011010011) && ({row_reg, col_reg}<16'b1001000011010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000011010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001000011010111) && ({row_reg, col_reg}<16'b1001000011011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000011011110) && ({row_reg, col_reg}<16'b1001000011100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001000011100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000011100010) && ({row_reg, col_reg}<16'b1001000011100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001000011100101) && ({row_reg, col_reg}<16'b1001000011100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000011100111) && ({row_reg, col_reg}<16'b1001000011101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001000011101001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001000011101010) && ({row_reg, col_reg}<16'b1001000011101100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==16'b1001000011101100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=16'b1001000011101101) && ({row_reg, col_reg}<16'b1001000011101111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001000011101111) && ({row_reg, col_reg}<16'b1001000011110100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001000011110100) && ({row_reg, col_reg}<16'b1001000011110110)) color_data = 12'b010000100001;

		if(({row_reg, col_reg}>=16'b1001000011110110) && ({row_reg, col_reg}<16'b1001000100000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001000100000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000100000001) && ({row_reg, col_reg}<16'b1001000100000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000100000011) && ({row_reg, col_reg}<16'b1001000100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001000100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000100000111) && ({row_reg, col_reg}<16'b1001000100001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001000100001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000100001010) && ({row_reg, col_reg}<16'b1001000100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000100001100) && ({row_reg, col_reg}<16'b1001000100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000100010001) && ({row_reg, col_reg}<16'b1001000100010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001000100010100) && ({row_reg, col_reg}<16'b1001000101100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001000101100100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001000101100101) && ({row_reg, col_reg}<16'b1001000101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001000101101001) && ({row_reg, col_reg}<16'b1001000101101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001000101101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000101101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000101101110) && ({row_reg, col_reg}<16'b1001000101111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000101111010) && ({row_reg, col_reg}<16'b1001000101111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001000101111100) && ({row_reg, col_reg}<16'b1001000101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001000101111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001000101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000110000000) && ({row_reg, col_reg}<16'b1001000110000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000110000100) && ({row_reg, col_reg}<16'b1001000110000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000110000110) && ({row_reg, col_reg}<16'b1001000110001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000110001000) && ({row_reg, col_reg}<16'b1001000110001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000110001010) && ({row_reg, col_reg}<16'b1001000110001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001000110001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000110001101) && ({row_reg, col_reg}<16'b1001000110010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001000110010011) && ({row_reg, col_reg}<16'b1001000110010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000110010110) && ({row_reg, col_reg}<16'b1001000110011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000110011000) && ({row_reg, col_reg}<16'b1001000110011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000110011010) && ({row_reg, col_reg}<16'b1001000110100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000110100010) && ({row_reg, col_reg}<16'b1001000110100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000110100110) && ({row_reg, col_reg}<16'b1001000110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000110110000) && ({row_reg, col_reg}<16'b1001000110110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001000110110011) && ({row_reg, col_reg}<16'b1001000110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000110110101) && ({row_reg, col_reg}<16'b1001000110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001000110111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001000110111111) && ({row_reg, col_reg}<16'b1001000111000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001000111000001) && ({row_reg, col_reg}<16'b1001000111000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000111000111) && ({row_reg, col_reg}<16'b1001000111001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001000111001101) && ({row_reg, col_reg}<16'b1001000111010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000111010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001000111010110) && ({row_reg, col_reg}<16'b1001000111011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000111011000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001000111011001) && ({row_reg, col_reg}<16'b1001000111011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001000111011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001000111011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000111011111) && ({row_reg, col_reg}<16'b1001000111101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001000111101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001000111101001) && ({row_reg, col_reg}<16'b1001000111101101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001000111101101) && ({row_reg, col_reg}<16'b1001000111110000)) color_data = 12'b010000100001;

		if(({row_reg, col_reg}>=16'b1001000111110000) && ({row_reg, col_reg}<16'b1001001000000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001001000000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001000000001) && ({row_reg, col_reg}<16'b1001001000000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001000000011) && ({row_reg, col_reg}<16'b1001001000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001000000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001000000110) && ({row_reg, col_reg}<16'b1001001000001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001000001001) && ({row_reg, col_reg}<16'b1001001000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001000001100) && ({row_reg, col_reg}<16'b1001001000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001000010001) && ({row_reg, col_reg}<16'b1001001000010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001001000010011) && ({row_reg, col_reg}<16'b1001001001101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001001001101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001001001101010) && ({row_reg, col_reg}<16'b1001001001101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001001101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001001001101101) && ({row_reg, col_reg}<16'b1001001001101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001001101111) && ({row_reg, col_reg}<16'b1001001001111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001001111010) && ({row_reg, col_reg}<16'b1001001001111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001001001111100) && ({row_reg, col_reg}<16'b1001001001111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001001001111111) && ({row_reg, col_reg}<16'b1001001010000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001001010000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001001010000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001010000110) && ({row_reg, col_reg}<16'b1001001010001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001010001000) && ({row_reg, col_reg}<16'b1001001010001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001001010001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001010001011) && ({row_reg, col_reg}<16'b1001001010001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001010001110) && ({row_reg, col_reg}<16'b1001001010010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001001010010010) && ({row_reg, col_reg}<16'b1001001010010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001010010101) && ({row_reg, col_reg}<16'b1001001010010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001010010111) && ({row_reg, col_reg}<16'b1001001010011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001010011010) && ({row_reg, col_reg}<16'b1001001010100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001010100010) && ({row_reg, col_reg}<16'b1001001010100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001010100110) && ({row_reg, col_reg}<16'b1001001010110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001010110001) && ({row_reg, col_reg}<16'b1001001010110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001010110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001010110101) && ({row_reg, col_reg}<16'b1001001010111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001010111111) && ({row_reg, col_reg}<16'b1001001011000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001001011000001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1001001011000010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001011000011) && ({row_reg, col_reg}<16'b1001001011000110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001001011000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001011000111) && ({row_reg, col_reg}<16'b1001001011001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001001011001100) && ({row_reg, col_reg}<16'b1001001011010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001011010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001001011010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001011010010) && ({row_reg, col_reg}<16'b1001001011010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001001011010100) && ({row_reg, col_reg}<16'b1001001011011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001011011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001001011011110) && ({row_reg, col_reg}<16'b1001001011100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001011100000) && ({row_reg, col_reg}<16'b1001001011100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001001011100110) && ({row_reg, col_reg}<16'b1001001011101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001011101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001001011101001) && ({row_reg, col_reg}<16'b1001001011101011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001011101011) && ({row_reg, col_reg}<16'b1001001011101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001001011101111) && ({row_reg, col_reg}<16'b1001001011110001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001001011110001) && ({row_reg, col_reg}<16'b1001001011111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001001011111010)) color_data = 12'b010000100001;

		if(({row_reg, col_reg}>=16'b1001001011111011) && ({row_reg, col_reg}<16'b1001001100000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001001100000000) && ({row_reg, col_reg}<16'b1001001100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001100000101) && ({row_reg, col_reg}<16'b1001001100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001100001100) && ({row_reg, col_reg}<16'b1001001100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001001100010010) && ({row_reg, col_reg}<16'b1001001101100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001001101100110) && ({row_reg, col_reg}<16'b1001001101101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001001101101001) && ({row_reg, col_reg}<16'b1001001101101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001001101101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001001101101101) && ({row_reg, col_reg}<16'b1001001101111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001101111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001001101111100) && ({row_reg, col_reg}<16'b1001001101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001001101111110) && ({row_reg, col_reg}<16'b1001001110000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001001110000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001001110000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001001110000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001110000110) && ({row_reg, col_reg}<16'b1001001110001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001001110001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001001110001010) && ({row_reg, col_reg}<16'b1001001110001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001110001111) && ({row_reg, col_reg}<16'b1001001110010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001001110010001) && ({row_reg, col_reg}<16'b1001001110010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001110010100) && ({row_reg, col_reg}<16'b1001001110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001110010111) && ({row_reg, col_reg}<16'b1001001110011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001110011101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001001110011110) && ({row_reg, col_reg}<16'b1001001110100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001110100011) && ({row_reg, col_reg}<16'b1001001110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001110101101) && ({row_reg, col_reg}<16'b1001001110110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001110110010) && ({row_reg, col_reg}<16'b1001001110111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001110111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001001110111100) && ({row_reg, col_reg}<16'b1001001111000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001001111000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001001111000010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001001111000011) && ({row_reg, col_reg}<16'b1001001111000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001111000110) && ({row_reg, col_reg}<16'b1001001111001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001001111001000) && ({row_reg, col_reg}<16'b1001001111001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001001111001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001001111001011)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==16'b1001001111001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001001111001101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001001111001110) && ({row_reg, col_reg}<16'b1001001111010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001111010000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001001111010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001001111010010)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==16'b1001001111010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001001111010100) && ({row_reg, col_reg}<16'b1001001111010111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001111010111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001001111011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001001111011001) && ({row_reg, col_reg}<16'b1001001111011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001001111011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001001111011100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001001111011101) && ({row_reg, col_reg}<16'b1001001111011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001111011111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001001111100000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001001111100001) && ({row_reg, col_reg}<16'b1001001111100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001001111100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001001111100110) && ({row_reg, col_reg}<16'b1001001111101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001001111101001) && ({row_reg, col_reg}<16'b1001001111101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001001111101011) && ({row_reg, col_reg}<16'b1001001111101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001001111101101) && ({row_reg, col_reg}<16'b1001001111101111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001001111101111) && ({row_reg, col_reg}<16'b1001001111110010)) color_data = 12'b010000110001;

		if(({row_reg, col_reg}>=16'b1001001111110010) && ({row_reg, col_reg}<16'b1001010000000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001010000000000) && ({row_reg, col_reg}<16'b1001010000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010000000101) && ({row_reg, col_reg}<16'b1001010000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010000001100) && ({row_reg, col_reg}<16'b1001010000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010000010001) && ({row_reg, col_reg}<16'b1001010001100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001010001100100) && ({row_reg, col_reg}<16'b1001010001100110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001010001100110) && ({row_reg, col_reg}<16'b1001010001101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010001101001) && ({row_reg, col_reg}<16'b1001010001101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010001101100) && ({row_reg, col_reg}<16'b1001010001101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001010001101110) && ({row_reg, col_reg}<16'b1001010001110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001010001110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001010001110100) && ({row_reg, col_reg}<16'b1001010001111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010001111001) && ({row_reg, col_reg}<16'b1001010001111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001010001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010001111110) && ({row_reg, col_reg}<16'b1001010010000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010010000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010010000100) && ({row_reg, col_reg}<16'b1001010010000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010010000110) && ({row_reg, col_reg}<16'b1001010010001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010010001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010010010000) && ({row_reg, col_reg}<16'b1001010010010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010010010010) && ({row_reg, col_reg}<16'b1001010010010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010010010111) && ({row_reg, col_reg}<16'b1001010010011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010010011010) && ({row_reg, col_reg}<16'b1001010010011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010010011100) && ({row_reg, col_reg}<16'b1001010010011110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010010011110) && ({row_reg, col_reg}<16'b1001010010100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010010100000) && ({row_reg, col_reg}<16'b1001010010100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001010010100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010010100011) && ({row_reg, col_reg}<16'b1001010010100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010010100101) && ({row_reg, col_reg}<16'b1001010010101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010010101101) && ({row_reg, col_reg}<16'b1001010010110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010010110011) && ({row_reg, col_reg}<16'b1001010010110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010010110101) && ({row_reg, col_reg}<16'b1001010010111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010010111001) && ({row_reg, col_reg}<16'b1001010011000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010011000010) && ({row_reg, col_reg}<16'b1001010011000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010011000100) && ({row_reg, col_reg}<16'b1001010011000111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001010011000111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010011001000) && ({row_reg, col_reg}<16'b1001010011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010011001010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001010011001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001010011001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010011001101) && ({row_reg, col_reg}<16'b1001010011010001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001010011010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010011010010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001010011010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010011010100) && ({row_reg, col_reg}<16'b1001010011011000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001010011011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010011011001) && ({row_reg, col_reg}<16'b1001010011011011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010011011011) && ({row_reg, col_reg}<16'b1001010011011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010011011101) && ({row_reg, col_reg}<16'b1001010011011111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001010011011111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010011100000) && ({row_reg, col_reg}<16'b1001010011100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010011100110) && ({row_reg, col_reg}<16'b1001010011101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010011101000) && ({row_reg, col_reg}<16'b1001010011101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010011101010) && ({row_reg, col_reg}<16'b1001010011101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010011101101) && ({row_reg, col_reg}<16'b1001010011101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010011101111) && ({row_reg, col_reg}<16'b1001010011110101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001010011110101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001010011110110) && ({row_reg, col_reg}<16'b1001010011111000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001010011111000) && ({row_reg, col_reg}<16'b1001010011111010)) color_data = 12'b010000100001;

		if(({row_reg, col_reg}>=16'b1001010011111010) && ({row_reg, col_reg}<16'b1001010100000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001010100000000) && ({row_reg, col_reg}<16'b1001010100000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010100000011) && ({row_reg, col_reg}<16'b1001010100000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001010100000101) && ({row_reg, col_reg}<16'b1001010100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010100001101) && ({row_reg, col_reg}<16'b1001010100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010100010001) && ({row_reg, col_reg}<16'b1001010101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001010101100011) && ({row_reg, col_reg}<16'b1001010101101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010101101000) && ({row_reg, col_reg}<16'b1001010101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010101101100) && ({row_reg, col_reg}<16'b1001010101101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001010101101110) && ({row_reg, col_reg}<16'b1001010101110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010101110010) && ({row_reg, col_reg}<16'b1001010101110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001010101110100) && ({row_reg, col_reg}<16'b1001010101111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010101111001) && ({row_reg, col_reg}<16'b1001010101111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001010101111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001010101111100) && ({row_reg, col_reg}<16'b1001010101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001010101111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001010110000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010110000001) && ({row_reg, col_reg}<16'b1001010110000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010110000110) && ({row_reg, col_reg}<16'b1001010110001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010110001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001010110001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001010110001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010110001101) && ({row_reg, col_reg}<16'b1001010110001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001010110001111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010110010000) && ({row_reg, col_reg}<16'b1001010110010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010110010010) && ({row_reg, col_reg}<16'b1001010110010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001010110010100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010110010101) && ({row_reg, col_reg}<16'b1001010110011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010110011101) && ({row_reg, col_reg}<16'b1001010110011111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010110011111) && ({row_reg, col_reg}<16'b1001010110100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001010110100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010110100101) && ({row_reg, col_reg}<16'b1001010110100111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001010110100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010110101000) && ({row_reg, col_reg}<16'b1001010110101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010110101101) && ({row_reg, col_reg}<16'b1001010110101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010110101111) && ({row_reg, col_reg}<16'b1001010110110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010110110101) && ({row_reg, col_reg}<16'b1001010110111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001010110111010) && ({row_reg, col_reg}<16'b1001010111000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010111000011) && ({row_reg, col_reg}<16'b1001010111000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010111000101) && ({row_reg, col_reg}<16'b1001010111001000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010111001000) && ({row_reg, col_reg}<16'b1001010111001100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010111001100) && ({row_reg, col_reg}<16'b1001010111010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001010111010101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001010111010110) && ({row_reg, col_reg}<16'b1001010111011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001010111011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001010111011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010111011110) && ({row_reg, col_reg}<16'b1001010111100000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001010111100000) && ({row_reg, col_reg}<16'b1001010111100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010111100011) && ({row_reg, col_reg}<16'b1001010111100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010111100101) && ({row_reg, col_reg}<16'b1001010111100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010111100111) && ({row_reg, col_reg}<16'b1001010111101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001010111101001) && ({row_reg, col_reg}<16'b1001010111101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001010111101011) && ({row_reg, col_reg}<16'b1001010111101111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001010111101111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001010111110000) && ({row_reg, col_reg}<16'b1001010111110110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001010111110110) && ({row_reg, col_reg}<16'b1001010111111100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001010111111100) && ({row_reg, col_reg}<16'b1001010111111111)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}==16'b1001010111111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011000000000) && ({row_reg, col_reg}<16'b1001011000000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001011000000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001011000000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011000000101) && ({row_reg, col_reg}<16'b1001011000001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011000001110) && ({row_reg, col_reg}<16'b1001011000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011000010001) && ({row_reg, col_reg}<16'b1001011001100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001011001100010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001011001100011) && ({row_reg, col_reg}<16'b1001011001101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011001101001) && ({row_reg, col_reg}<16'b1001011001101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011001101100) && ({row_reg, col_reg}<16'b1001011001101110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001011001101110) && ({row_reg, col_reg}<16'b1001011001110010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011001110010) && ({row_reg, col_reg}<16'b1001011001110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001011001110101) && ({row_reg, col_reg}<16'b1001011001110111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011001110111) && ({row_reg, col_reg}<16'b1001011001111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001011001111001) && ({row_reg, col_reg}<16'b1001011001111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001011001111011) && ({row_reg, col_reg}<16'b1001011001111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011001111101) && ({row_reg, col_reg}<16'b1001011010000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011010000010) && ({row_reg, col_reg}<16'b1001011010000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011010000110) && ({row_reg, col_reg}<16'b1001011010001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011010001010) && ({row_reg, col_reg}<16'b1001011010001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001011010001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011010001111) && ({row_reg, col_reg}<16'b1001011010010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001011010010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011010010011) && ({row_reg, col_reg}<16'b1001011010010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011010010101) && ({row_reg, col_reg}<16'b1001011010011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011010011101) && ({row_reg, col_reg}<16'b1001011010100100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011010100100) && ({row_reg, col_reg}<16'b1001011010101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011010101000) && ({row_reg, col_reg}<16'b1001011010101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011010101100) && ({row_reg, col_reg}<16'b1001011010101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011010101110) && ({row_reg, col_reg}<16'b1001011010110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011010110011) && ({row_reg, col_reg}<16'b1001011010110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011010110101) && ({row_reg, col_reg}<16'b1001011010111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011010111010) && ({row_reg, col_reg}<16'b1001011011000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011011000100) && ({row_reg, col_reg}<16'b1001011011000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001011011000110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001011011000111) && ({row_reg, col_reg}<16'b1001011011001001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011011001001) && ({row_reg, col_reg}<16'b1001011011001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001011011001011) && ({row_reg, col_reg}<16'b1001011011011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001011011011001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001011011011010) && ({row_reg, col_reg}<16'b1001011011011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011011011100) && ({row_reg, col_reg}<16'b1001011011011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001011011011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001011011011111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001011011100000) && ({row_reg, col_reg}<16'b1001011011100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011011100011) && ({row_reg, col_reg}<16'b1001011011100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011011100101) && ({row_reg, col_reg}<16'b1001011011100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011011100111) && ({row_reg, col_reg}<16'b1001011011101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011011101011) && ({row_reg, col_reg}<16'b1001011011110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001011011110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011011110001) && ({row_reg, col_reg}<16'b1001011011110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011011110011) && ({row_reg, col_reg}<16'b1001011011110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001011011110111) && ({row_reg, col_reg}<16'b1001011011111001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=16'b1001011011111001) && ({row_reg, col_reg}<16'b1001011011111110)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}>=16'b1001011011111110) && ({row_reg, col_reg}<16'b1001011100000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011100000000) && ({row_reg, col_reg}<16'b1001011100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011100000110) && ({row_reg, col_reg}<16'b1001011100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001011100001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011100001100) && ({row_reg, col_reg}<16'b1001011100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011100001111) && ({row_reg, col_reg}<16'b1001011100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001011100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001011100010010) && ({row_reg, col_reg}<16'b1001011101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001011101100011) && ({row_reg, col_reg}<16'b1001011101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011101101010) && ({row_reg, col_reg}<16'b1001011101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001011101101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001011101101101) && ({row_reg, col_reg}<16'b1001011101110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011101110011) && ({row_reg, col_reg}<16'b1001011101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001011101110110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011101110111) && ({row_reg, col_reg}<16'b1001011101111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001011101111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011101111010) && ({row_reg, col_reg}<16'b1001011101111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011101111110) && ({row_reg, col_reg}<16'b1001011110000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011110000000) && ({row_reg, col_reg}<16'b1001011110001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011110001110) && ({row_reg, col_reg}<16'b1001011110010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001011110010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011110010001) && ({row_reg, col_reg}<16'b1001011110010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011110010110) && ({row_reg, col_reg}<16'b1001011110011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011110011011) && ({row_reg, col_reg}<16'b1001011110100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011110100001) && ({row_reg, col_reg}<16'b1001011110101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011110101110) && ({row_reg, col_reg}<16'b1001011110110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011110110100) && ({row_reg, col_reg}<16'b1001011110111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011110111101) && ({row_reg, col_reg}<16'b1001011111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011111000101) && ({row_reg, col_reg}<16'b1001011111000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011111000111) && ({row_reg, col_reg}<16'b1001011111001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001011111001001) && ({row_reg, col_reg}<16'b1001011111010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001011111010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001011111010010) && ({row_reg, col_reg}<16'b1001011111011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001011111011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001011111011001) && ({row_reg, col_reg}<16'b1001011111011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011111011100) && ({row_reg, col_reg}<16'b1001011111011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001011111011110) && ({row_reg, col_reg}<16'b1001011111100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001011111100000) && ({row_reg, col_reg}<16'b1001011111100111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011111100111) && ({row_reg, col_reg}<16'b1001011111101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001011111101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001011111101010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011111101011) && ({row_reg, col_reg}<16'b1001011111101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001011111101111) && ({row_reg, col_reg}<16'b1001011111110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001011111110011) && ({row_reg, col_reg}<16'b1001011111110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011111110101) && ({row_reg, col_reg}<16'b1001011111111100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001011111111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001011111111101) && ({row_reg, col_reg}<16'b1001011111111111)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}==16'b1001011111111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100000000000) && ({row_reg, col_reg}<16'b1001100000000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100000000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100000000110) && ({row_reg, col_reg}<16'b1001100000001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100000001111) && ({row_reg, col_reg}<16'b1001100000010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001100000010010) && ({row_reg, col_reg}<16'b1001100001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001100001100011) && ({row_reg, col_reg}<16'b1001100001101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100001101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001100001101101) && ({row_reg, col_reg}<16'b1001100001110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100001110011) && ({row_reg, col_reg}<16'b1001100001111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001100001111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100001111001) && ({row_reg, col_reg}<16'b1001100001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100001111011) && ({row_reg, col_reg}<16'b1001100010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100010000010) && ({row_reg, col_reg}<16'b1001100010001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100010001100) && ({row_reg, col_reg}<16'b1001100010010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100010010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100010010001) && ({row_reg, col_reg}<16'b1001100010011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100010011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100010011011) && ({row_reg, col_reg}<16'b1001100010100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100010100110) && ({row_reg, col_reg}<16'b1001100010101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100010101011) && ({row_reg, col_reg}<16'b1001100010110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100010110100) && ({row_reg, col_reg}<16'b1001100010111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100010111111) && ({row_reg, col_reg}<16'b1001100011000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100011000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100011001000) && ({row_reg, col_reg}<16'b1001100011001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001100011001010) && ({row_reg, col_reg}<16'b1001100011010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100011010010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001100011010011) && ({row_reg, col_reg}<16'b1001100011011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100011011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001100011011001) && ({row_reg, col_reg}<16'b1001100011011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100011011110) && ({row_reg, col_reg}<16'b1001100011100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001100011100000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100011100001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001100011100010) && ({row_reg, col_reg}<16'b1001100011100110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100011100110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1001100011100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100011101000) && ({row_reg, col_reg}<16'b1001100011101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100011101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001100011101011) && ({row_reg, col_reg}<16'b1001100011110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001100011110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001100011110110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100011110111) && ({row_reg, col_reg}<16'b1001100011111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001100011111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100011111011) && ({row_reg, col_reg}<16'b1001100011111111)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}==16'b1001100011111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100100000000) && ({row_reg, col_reg}<16'b1001100100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100100000101) && ({row_reg, col_reg}<16'b1001100100000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100100000111) && ({row_reg, col_reg}<16'b1001100100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001100100001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100100001100) && ({row_reg, col_reg}<16'b1001100100001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100100001110) && ({row_reg, col_reg}<16'b1001100100010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001100100010010) && ({row_reg, col_reg}<16'b1001100101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001100101100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001100101100100) && ({row_reg, col_reg}<16'b1001100101101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100101101000) && ({row_reg, col_reg}<16'b1001100101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001100101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100101101011) && ({row_reg, col_reg}<16'b1001100101101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001100101101101) && ({row_reg, col_reg}<16'b1001100101110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100101110011) && ({row_reg, col_reg}<16'b1001100101110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001100101110110) && ({row_reg, col_reg}<16'b1001100101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100101111000) && ({row_reg, col_reg}<16'b1001100101111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001100101111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001100101111011) && ({row_reg, col_reg}<16'b1001100101111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100101111101) && ({row_reg, col_reg}<16'b1001100110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100110000010) && ({row_reg, col_reg}<16'b1001100110001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100110001011) && ({row_reg, col_reg}<16'b1001100110001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100110001101) && ({row_reg, col_reg}<16'b1001100110010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100110010110) && ({row_reg, col_reg}<16'b1001100110011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100110011101) && ({row_reg, col_reg}<16'b1001100110100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100110100110) && ({row_reg, col_reg}<16'b1001100110101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100110101011) && ({row_reg, col_reg}<16'b1001100110101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100110101111) && ({row_reg, col_reg}<16'b1001100110111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100110111110) && ({row_reg, col_reg}<16'b1001100111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001100111001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100111001010) && ({row_reg, col_reg}<16'b1001100111011000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100111011000) && ({row_reg, col_reg}<16'b1001100111011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001100111011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100111011101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001100111011110) && ({row_reg, col_reg}<16'b1001100111100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001100111100000) && ({row_reg, col_reg}<16'b1001100111100100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100111100100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001100111100101) && ({row_reg, col_reg}<16'b1001100111101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100111101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001100111101010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001100111101011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100111101100) && ({row_reg, col_reg}<16'b1001100111110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001100111110011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001100111110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001100111110101) && ({row_reg, col_reg}<16'b1001100111110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001100111110111) && ({row_reg, col_reg}<16'b1001100111111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001100111111010) && ({row_reg, col_reg}<16'b1001100111111111)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}==16'b1001100111111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101000000000) && ({row_reg, col_reg}<16'b1001101000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101000000110) && ({row_reg, col_reg}<16'b1001101000001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101000001010) && ({row_reg, col_reg}<16'b1001101000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101000001111) && ({row_reg, col_reg}<16'b1001101000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001101000010010) && ({row_reg, col_reg}<16'b1001101001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001101001100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001101001100100) && ({row_reg, col_reg}<16'b1001101001101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101001101000) && ({row_reg, col_reg}<16'b1001101001101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101001101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101001101011) && ({row_reg, col_reg}<16'b1001101001101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001101001101101) && ({row_reg, col_reg}<16'b1001101001110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101001110011) && ({row_reg, col_reg}<16'b1001101001110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001101001110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001101001110110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101001110111) && ({row_reg, col_reg}<16'b1001101001111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001101001111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101001111010) && ({row_reg, col_reg}<16'b1001101001111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001101001111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101010000000) && ({row_reg, col_reg}<16'b1001101010000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101010000011) && ({row_reg, col_reg}<16'b1001101010000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101010000101) && ({row_reg, col_reg}<16'b1001101010000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101010000111) && ({row_reg, col_reg}<16'b1001101010001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101010001011) && ({row_reg, col_reg}<16'b1001101010010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101010010011) && ({row_reg, col_reg}<16'b1001101010010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101010010101) && ({row_reg, col_reg}<16'b1001101010011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101010011101) && ({row_reg, col_reg}<16'b1001101010100110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101010100110) && ({row_reg, col_reg}<16'b1001101010101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101010101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101010101010) && ({row_reg, col_reg}<16'b1001101010101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101010101111) && ({row_reg, col_reg}<16'b1001101010110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101010110111) && ({row_reg, col_reg}<16'b1001101010111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101010111010) && ({row_reg, col_reg}<16'b1001101010111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101010111101) && ({row_reg, col_reg}<16'b1001101011000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101011000000) && ({row_reg, col_reg}<16'b1001101011000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101011000010) && ({row_reg, col_reg}<16'b1001101011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001101011001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101011001011) && ({row_reg, col_reg}<16'b1001101011001110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001101011001110) && ({row_reg, col_reg}<16'b1001101011011001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101011011001) && ({row_reg, col_reg}<16'b1001101011011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001101011011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101011011101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101011011110) && ({row_reg, col_reg}<16'b1001101011100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101011100000) && ({row_reg, col_reg}<16'b1001101011100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101011100101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001101011100110) && ({row_reg, col_reg}<16'b1001101011101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101011101000) && ({row_reg, col_reg}<16'b1001101011101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001101011101010) && ({row_reg, col_reg}<16'b1001101011101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101011101101) && ({row_reg, col_reg}<16'b1001101011101111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001101011101111) && ({row_reg, col_reg}<16'b1001101011110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101011110011) && ({row_reg, col_reg}<16'b1001101011111100)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}>=16'b1001101011111100) && ({row_reg, col_reg}<16'b1001101100000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101100000001) && ({row_reg, col_reg}<16'b1001101100000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101100000111) && ({row_reg, col_reg}<16'b1001101100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101100001001) && ({row_reg, col_reg}<16'b1001101100001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101100001101) && ({row_reg, col_reg}<16'b1001101100001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001101100001111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001101100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101100010001) && ({row_reg, col_reg}<16'b1001101101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001101101100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001101101100100) && ({row_reg, col_reg}<16'b1001101101101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101101101000) && ({row_reg, col_reg}<16'b1001101101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101101101011) && ({row_reg, col_reg}<16'b1001101101101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001101101101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001101101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101101101111) && ({row_reg, col_reg}<16'b1001101101110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101101110101) && ({row_reg, col_reg}<16'b1001101101110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001101101110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101101111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001101101111001) && ({row_reg, col_reg}<16'b1001101101111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001101101111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101110000000) && ({row_reg, col_reg}<16'b1001101110000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101110000011) && ({row_reg, col_reg}<16'b1001101110000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101110000101) && ({row_reg, col_reg}<16'b1001101110000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101110000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001101110001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101110001001) && ({row_reg, col_reg}<16'b1001101110001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101110001101) && ({row_reg, col_reg}<16'b1001101110010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101110010010) && ({row_reg, col_reg}<16'b1001101110010110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101110010110) && ({row_reg, col_reg}<16'b1001101110011011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101110011011) && ({row_reg, col_reg}<16'b1001101110011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101110011110) && ({row_reg, col_reg}<16'b1001101110100001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001101110100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101110100010) && ({row_reg, col_reg}<16'b1001101110100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001101110100101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101110100110) && ({row_reg, col_reg}<16'b1001101110101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101110101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101110101010) && ({row_reg, col_reg}<16'b1001101110101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101110101100) && ({row_reg, col_reg}<16'b1001101110101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101110101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101110101111) && ({row_reg, col_reg}<16'b1001101110110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101110110111) && ({row_reg, col_reg}<16'b1001101110111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001101110111010) && ({row_reg, col_reg}<16'b1001101110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001101110111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101110111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101111000000) && ({row_reg, col_reg}<16'b1001101111000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101111000010) && ({row_reg, col_reg}<16'b1001101111001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101111001100) && ({row_reg, col_reg}<16'b1001101111001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001101111001110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001101111001111) && ({row_reg, col_reg}<16'b1001101111010001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101111010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001101111010010) && ({row_reg, col_reg}<16'b1001101111011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101111011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001101111011100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001101111011101) && ({row_reg, col_reg}<16'b1001101111011111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101111011111) && ({row_reg, col_reg}<16'b1001101111100001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001101111100001) && ({row_reg, col_reg}<16'b1001101111101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101111101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001101111101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101111101010) && ({row_reg, col_reg}<16'b1001101111101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001101111101100) && ({row_reg, col_reg}<16'b1001101111110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001101111110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001101111110001) && ({row_reg, col_reg}<16'b1001101111110011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001101111110011) && ({row_reg, col_reg}<16'b1001101111111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001101111111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001101111111001) && ({row_reg, col_reg}<16'b1001101111111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001101111111011) && ({row_reg, col_reg}<16'b1001101111111111)) color_data = 12'b001000100001;

		if(({row_reg, col_reg}==16'b1001101111111111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1001110000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110000000001) && ({row_reg, col_reg}<16'b1001110000000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110000000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110000001000) && ({row_reg, col_reg}<16'b1001110000001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110000001011) && ({row_reg, col_reg}<16'b1001110000001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110000001101) && ({row_reg, col_reg}<16'b1001110000010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001110000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001110000010010) && ({row_reg, col_reg}<16'b1001110001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001110001100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001110001100100) && ({row_reg, col_reg}<16'b1001110001101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110001101000) && ({row_reg, col_reg}<16'b1001110001101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110001101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110001101011) && ({row_reg, col_reg}<16'b1001110001101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001110001101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110001101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110001101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110001110000) && ({row_reg, col_reg}<16'b1001110001110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001110001110010) && ({row_reg, col_reg}<16'b1001110001110100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110001110100) && ({row_reg, col_reg}<16'b1001110001110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001110001110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==16'b1001110001111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110001111001) && ({row_reg, col_reg}<16'b1001110010000000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110010000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110010000001) && ({row_reg, col_reg}<16'b1001110010000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110010000011) && ({row_reg, col_reg}<16'b1001110010000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110010000110) && ({row_reg, col_reg}<16'b1001110010001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110010001101) && ({row_reg, col_reg}<16'b1001110010010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110010010010) && ({row_reg, col_reg}<16'b1001110010010101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110010010101) && ({row_reg, col_reg}<16'b1001110010011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110010011010) && ({row_reg, col_reg}<16'b1001110010011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110010011110) && ({row_reg, col_reg}<16'b1001110010100000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001110010100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110010100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110010100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110010100011) && ({row_reg, col_reg}<16'b1001110010100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110010100101) && ({row_reg, col_reg}<16'b1001110010101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110010101110) && ({row_reg, col_reg}<16'b1001110010111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110010111010) && ({row_reg, col_reg}<16'b1001110010111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110010111101) && ({row_reg, col_reg}<16'b1001110010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110010111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110011000000) && ({row_reg, col_reg}<16'b1001110011000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110011000010) && ({row_reg, col_reg}<16'b1001110011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110011001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001110011001111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1001110011010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110011010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001110011010010) && ({row_reg, col_reg}<16'b1001110011010101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110011010101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001110011010110) && ({row_reg, col_reg}<16'b1001110011011011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110011011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001110011011100) && ({row_reg, col_reg}<16'b1001110011011110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001110011011110) && ({row_reg, col_reg}<16'b1001110011100000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001110011100000) && ({row_reg, col_reg}<16'b1001110011100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110011100011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001110011100100) && ({row_reg, col_reg}<16'b1001110011101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110011101010) && ({row_reg, col_reg}<16'b1001110011101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001110011101100) && ({row_reg, col_reg}<16'b1001110011110000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110011110000) && ({row_reg, col_reg}<16'b1001110011110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001110011110010) && ({row_reg, col_reg}<16'b1001110011110111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110011110111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001110011111000) && ({row_reg, col_reg}<16'b1001110011111010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110011111010) && ({row_reg, col_reg}<16'b1001110011111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110011111100) && ({row_reg, col_reg}<16'b1001110011111110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001110011111110)) color_data = 12'b001000100001;

		if(({row_reg, col_reg}==16'b1001110011111111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=16'b1001110100000000) && ({row_reg, col_reg}<16'b1001110100000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110100000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110100000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110100001000) && ({row_reg, col_reg}<16'b1001110100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001110100001100) && ({row_reg, col_reg}<16'b1001110100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110100001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001110100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001110100010010) && ({row_reg, col_reg}<16'b1001110101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001110101100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001110101100100) && ({row_reg, col_reg}<16'b1001110101101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110101101000) && ({row_reg, col_reg}<16'b1001110101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110101101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==16'b1001110101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001110101101101) && ({row_reg, col_reg}<16'b1001110101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110101110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001110101110001) && ({row_reg, col_reg}<16'b1001110101110011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110101110011) && ({row_reg, col_reg}<16'b1001110101111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110101111001) && ({row_reg, col_reg}<16'b1001110110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110110000010) && ({row_reg, col_reg}<16'b1001110110000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110110000110) && ({row_reg, col_reg}<16'b1001110110001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110110001100) && ({row_reg, col_reg}<16'b1001110110011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110110011010) && ({row_reg, col_reg}<16'b1001110110011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110110011101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001110110011110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001110110011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110110100000) && ({row_reg, col_reg}<16'b1001110110100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110110100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110110100011) && ({row_reg, col_reg}<16'b1001110110100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110110100101) && ({row_reg, col_reg}<16'b1001110110101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110110101100) && ({row_reg, col_reg}<16'b1001110110111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001110110111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110110111100) && ({row_reg, col_reg}<16'b1001110110111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001110110111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110111000000) && ({row_reg, col_reg}<16'b1001110111000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110111000011) && ({row_reg, col_reg}<16'b1001110111001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001110111001110) && ({row_reg, col_reg}<16'b1001110111010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110111010000) && ({row_reg, col_reg}<16'b1001110111010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110111010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001110111010100) && ({row_reg, col_reg}<16'b1001110111010110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110111010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001110111010111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b1001110111011000) && ({row_reg, col_reg}<16'b1001110111011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001110111011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110111011011) && ({row_reg, col_reg}<16'b1001110111011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001110111011101) && ({row_reg, col_reg}<16'b1001110111100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110111100011) && ({row_reg, col_reg}<16'b1001110111100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001110111100101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110111100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001110111100111) && ({row_reg, col_reg}<16'b1001110111101001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110111101001) && ({row_reg, col_reg}<16'b1001110111101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001110111101011) && ({row_reg, col_reg}<16'b1001110111101101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110111101101) && ({row_reg, col_reg}<16'b1001110111101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001110111101111) && ({row_reg, col_reg}<16'b1001110111110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110111110101) && ({row_reg, col_reg}<16'b1001110111110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001110111110111) && ({row_reg, col_reg}<16'b1001110111111001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001110111111001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001110111111010) && ({row_reg, col_reg}<16'b1001110111111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001110111111100) && ({row_reg, col_reg}<16'b1001110111111111)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}==16'b1001110111111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111000000000) && ({row_reg, col_reg}<16'b1001111000000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111000000010) && ({row_reg, col_reg}<16'b1001111000000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001111000000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111000000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001111000000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111000000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001111000001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111000001001) && ({row_reg, col_reg}<16'b1001111000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111000001100) && ({row_reg, col_reg}<16'b1001111000001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111000001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001111000010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111000010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001111000010010) && ({row_reg, col_reg}<16'b1001111001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001111001100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001111001100100) && ({row_reg, col_reg}<16'b1001111001101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111001101000) && ({row_reg, col_reg}<16'b1001111001101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001111001101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111001101011) && ({row_reg, col_reg}<16'b1001111001101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001111001101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001111001101110) && ({row_reg, col_reg}<16'b1001111001110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111001110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001111001110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001111001110011) && ({row_reg, col_reg}<16'b1001111001110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001111001110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111001110110) && ({row_reg, col_reg}<16'b1001111001111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111001111000) && ({row_reg, col_reg}<16'b1001111001111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111001111110) && ({row_reg, col_reg}<16'b1001111010000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111010000000) && ({row_reg, col_reg}<16'b1001111010000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111010000010) && ({row_reg, col_reg}<16'b1001111010000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111010000110) && ({row_reg, col_reg}<16'b1001111010001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111010001000) && ({row_reg, col_reg}<16'b1001111010001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001111010001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111010001011) && ({row_reg, col_reg}<16'b1001111010011110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001111010011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111010011111) && ({row_reg, col_reg}<16'b1001111010100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001111010100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111010100011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111010100100) && ({row_reg, col_reg}<16'b1001111010101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111010101010) && ({row_reg, col_reg}<16'b1001111010101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111010101101) && ({row_reg, col_reg}<16'b1001111010111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001111010111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111010111100) && ({row_reg, col_reg}<16'b1001111010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001111010111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111011000000) && ({row_reg, col_reg}<16'b1001111011000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111011000100) && ({row_reg, col_reg}<16'b1001111011010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111011010000) && ({row_reg, col_reg}<16'b1001111011010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001111011010010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111011010011) && ({row_reg, col_reg}<16'b1001111011010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001111011010110) && ({row_reg, col_reg}<16'b1001111011011000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b1001111011011000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==16'b1001111011011001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001111011011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111011011011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b1001111011011100) && ({row_reg, col_reg}<16'b1001111011011110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b1001111011011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001111011011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111011100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001111011100001) && ({row_reg, col_reg}<16'b1001111011100011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111011100011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==16'b1001111011100100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001111011100101) && ({row_reg, col_reg}<16'b1001111011101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111011101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001111011101001)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==16'b1001111011101010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001111011101011) && ({row_reg, col_reg}<16'b1001111011110001)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111011110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001111011110010) && ({row_reg, col_reg}<16'b1001111011110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111011110101) && ({row_reg, col_reg}<16'b1001111011110111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001111011110111) && ({row_reg, col_reg}<16'b1001111011111100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111011111100) && ({row_reg, col_reg}<16'b1001111011111111)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}==16'b1001111011111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111100000000) && ({row_reg, col_reg}<16'b1001111100000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111100000110) && ({row_reg, col_reg}<16'b1001111100001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111100001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111100001001) && ({row_reg, col_reg}<16'b1001111100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111100001100) && ({row_reg, col_reg}<16'b1001111100001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111100001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001111100010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001111100010010) && ({row_reg, col_reg}<16'b1001111101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==16'b1001111101100011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001111101100100) && ({row_reg, col_reg}<16'b1001111101101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==16'b1001111101101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=16'b1001111101101011) && ({row_reg, col_reg}<16'b1001111101101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001111101101110) && ({row_reg, col_reg}<16'b1001111101110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111101110000) && ({row_reg, col_reg}<16'b1001111101110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001111101110010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=16'b1001111101110011) && ({row_reg, col_reg}<16'b1001111101110101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001111101110101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111101110110) && ({row_reg, col_reg}<16'b1001111101111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111101111000) && ({row_reg, col_reg}<16'b1001111110000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111110000010) && ({row_reg, col_reg}<16'b1001111110000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001111110000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111110000111) && ({row_reg, col_reg}<16'b1001111110001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111110001001) && ({row_reg, col_reg}<16'b1001111110001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111110001110) && ({row_reg, col_reg}<16'b1001111110010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111110010000) && ({row_reg, col_reg}<16'b1001111110010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111110010011) && ({row_reg, col_reg}<16'b1001111110011111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111110011111) && ({row_reg, col_reg}<16'b1001111110100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111110100010) && ({row_reg, col_reg}<16'b1001111110100101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111110100101) && ({row_reg, col_reg}<16'b1001111110101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111110101000) && ({row_reg, col_reg}<16'b1001111110101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=16'b1001111110101010) && ({row_reg, col_reg}<16'b1001111110101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111110101100) && ({row_reg, col_reg}<16'b1001111110111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001111110111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111110111100) && ({row_reg, col_reg}<16'b1001111110111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==16'b1001111110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111110111111) && ({row_reg, col_reg}<16'b1001111111000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=16'b1001111111000101) && ({row_reg, col_reg}<16'b1001111111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=16'b1001111111010001) && ({row_reg, col_reg}<16'b1001111111010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==16'b1001111111010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111111010100) && ({row_reg, col_reg}<16'b1001111111010110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=16'b1001111111010110) && ({row_reg, col_reg}<16'b1001111111011000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b1001111111011000) && ({row_reg, col_reg}<16'b1001111111011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001111111011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111111011011) && ({row_reg, col_reg}<16'b1001111111011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001111111011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111111100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001111111100001) && ({row_reg, col_reg}<16'b1001111111101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==16'b1001111111101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==16'b1001111111101001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=16'b1001111111101010) && ({row_reg, col_reg}<16'b1001111111101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==16'b1001111111101100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111111101101) && ({row_reg, col_reg}<16'b1001111111110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=16'b1001111111110000) && ({row_reg, col_reg}<16'b1001111111111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=16'b1001111111111010) && ({row_reg, col_reg}<16'b1001111111111100)) color_data = 12'b001000100000;

		if(({row_reg, col_reg}>=16'b1001111111111100) && ({row_reg, col_reg}<=16'b1001111111111111)) color_data = 12'b001100100001;
	end
endmodule