module shoot2_rom
	(
		input wire clk,
		input wire [6:0] row,
		input wire [6:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [6:0] row_reg;
	reg [6:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin
		if(({row_reg, col_reg}>=14'b00000000000000) && ({row_reg, col_reg}<14'b00000000110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00000000110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00000000110011) && ({row_reg, col_reg}<14'b00000000110101)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=14'b00000000110101) && ({row_reg, col_reg}<14'b00000010110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00000010110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00000010110010) && ({row_reg, col_reg}<14'b00000010110101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00000010110101) && ({row_reg, col_reg}<14'b00000010111000)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=14'b00000010111000) && ({row_reg, col_reg}<14'b00000100110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00000100110001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00000100110010) && ({row_reg, col_reg}<14'b00000100110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00000100110110) && ({row_reg, col_reg}<14'b00000100111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00000100111000) && ({row_reg, col_reg}<14'b00000100111010)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=14'b00000100111010) && ({row_reg, col_reg}<14'b00000110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00000110110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00000110110001) && ({row_reg, col_reg}<14'b00000110111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00000110111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00000110111001) && ({row_reg, col_reg}<14'b00000110111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00000110111101)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00000110111110) && ({row_reg, col_reg}<14'b00001000110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00001000110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00001000110001) && ({row_reg, col_reg}<14'b00001000110011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00001000110011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00001000110100) && ({row_reg, col_reg}<14'b00001000111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00001000111000) && ({row_reg, col_reg}<14'b00001000111101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00001000111101) && ({row_reg, col_reg}<14'b00001001000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00001001000000)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00001001000001) && ({row_reg, col_reg}<14'b00001010101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00001010101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00001010110000) && ({row_reg, col_reg}<14'b00001010111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00001010111000) && ({row_reg, col_reg}<14'b00001010111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00001010111011) && ({row_reg, col_reg}<14'b00001010111101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00001010111101) && ({row_reg, col_reg}<14'b00001010111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00001010111111) && ({row_reg, col_reg}<14'b00001011000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00001011000001)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00001011000010) && ({row_reg, col_reg}<14'b00001100101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00001100101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00001100110000) && ({row_reg, col_reg}<14'b00001100110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00001100110111) && ({row_reg, col_reg}<14'b00001100111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00001100111001) && ({row_reg, col_reg}<14'b00001100111111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00001100111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00001101000000) && ({row_reg, col_reg}<14'b00001101000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00001101000010)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00001101000011) && ({row_reg, col_reg}<14'b00001110101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b00001110101111) && ({row_reg, col_reg}<14'b00001110110101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00001110110101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00001110110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00001110110111) && ({row_reg, col_reg}<14'b00001110111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00001110111001) && ({row_reg, col_reg}<14'b00001110111011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00001110111011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b00001110111100) && ({row_reg, col_reg}<14'b00001110111111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00001110111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00001111000000) && ({row_reg, col_reg}<14'b00001111000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00001111000010) && ({row_reg, col_reg}<14'b00001111000100)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00001111000100) && ({row_reg, col_reg}<14'b00010000101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00010000101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00010000101111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b00010000110000) && ({row_reg, col_reg}<14'b00010000110101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00010000110101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00010000110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00010000110111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00010000111000) && ({row_reg, col_reg}<14'b00010000111010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00010000111010) && ({row_reg, col_reg}<14'b00010000111110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00010000111110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00010000111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00010001000000) && ({row_reg, col_reg}<14'b00010001000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00010001000011)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00010001000100) && ({row_reg, col_reg}<14'b00010010101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00010010101110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00010010101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b00010010110000) && ({row_reg, col_reg}<14'b00010010110110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b00010010110110) && ({row_reg, col_reg}<14'b00010010111001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00010010111001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b00010010111010) && ({row_reg, col_reg}<14'b00010010111101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00010010111101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b00010010111110) && ({row_reg, col_reg}<14'b00010011000000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00010011000000) && ({row_reg, col_reg}<14'b00010011000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00010011000100)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00010011000101) && ({row_reg, col_reg}<14'b00010100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00010100101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00010100101110) && ({row_reg, col_reg}<14'b00010100110000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b00010100110000) && ({row_reg, col_reg}<14'b00010100110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00010100110101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00010100110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00010100110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00010100111000) && ({row_reg, col_reg}<14'b00010100111010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b00010100111010) && ({row_reg, col_reg}<14'b00010100111101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b00010100111101) && ({row_reg, col_reg}<14'b00010100111111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00010100111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00010101000000) && ({row_reg, col_reg}<14'b00010101000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00010101000100)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00010101000101) && ({row_reg, col_reg}<14'b00010110101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00010110101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00010110101110) && ({row_reg, col_reg}<14'b00010110110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00010110110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b00010110110001) && ({row_reg, col_reg}<14'b00010110110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00010110110101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b00010110110110) && ({row_reg, col_reg}<14'b00010110111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00010110111000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00010110111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b00010110111010) && ({row_reg, col_reg}<14'b00010110111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00010110111100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00010110111101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00010110111110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00010110111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00010111000000) && ({row_reg, col_reg}<14'b00010111000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00010111000100)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00010111000101) && ({row_reg, col_reg}<14'b00011000101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b00011000101101) && ({row_reg, col_reg}<14'b00011000101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00011000101111) && ({row_reg, col_reg}<14'b00011000110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00011000110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00011000110010) && ({row_reg, col_reg}<14'b00011000110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00011000110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b00011000110101) && ({row_reg, col_reg}<14'b00011000111000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00011000111000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b00011000111001) && ({row_reg, col_reg}<14'b00011000111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00011000111100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00011000111101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00011000111110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00011000111111) && ({row_reg, col_reg}<14'b00011001000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00011001000100) && ({row_reg, col_reg}<14'b00011001000110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00011001000110) && ({row_reg, col_reg}<14'b00011010101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b00011010101101) && ({row_reg, col_reg}<14'b00011010110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00011010110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00011010110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00011010110011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b00011010110100) && ({row_reg, col_reg}<14'b00011010110110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b00011010110110) && ({row_reg, col_reg}<14'b00011010111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b00011010111001) && ({row_reg, col_reg}<14'b00011010111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00011010111100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00011010111101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00011010111110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00011010111111) && ({row_reg, col_reg}<14'b00011011000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00011011000100) && ({row_reg, col_reg}<14'b00011011000110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00011011000110) && ({row_reg, col_reg}<14'b00011100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b00011100101100) && ({row_reg, col_reg}<14'b00011100110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00011100110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00011100110011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00011100110100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00011100110101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b00011100110110) && ({row_reg, col_reg}<14'b00011100111000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00011100111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00011100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b00011100111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b00011100111011) && ({row_reg, col_reg}<14'b00011100111101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00011100111101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00011100111110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00011100111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00011101000000) && ({row_reg, col_reg}<14'b00011101000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00011101000101)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00011101000110) && ({row_reg, col_reg}<14'b00011110101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b00011110101100) && ({row_reg, col_reg}<14'b00011110110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00011110110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00011110110011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00011110110100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00011110110101) && ({row_reg, col_reg}<14'b00011110110111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b00011110110111) && ({row_reg, col_reg}<14'b00011110111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b00011110111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b00011110111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b00011110111011) && ({row_reg, col_reg}<14'b00011110111101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00011110111101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00011110111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00011110111111) && ({row_reg, col_reg}<14'b00011111000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00011111000100) && ({row_reg, col_reg}<14'b00011111000110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00011111000110) && ({row_reg, col_reg}<14'b00100000101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b00100000101011) && ({row_reg, col_reg}<14'b00100000110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00100000110000) && ({row_reg, col_reg}<14'b00100000110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00100000110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00100000110100) && ({row_reg, col_reg}<14'b00100000111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00100000111000) && ({row_reg, col_reg}<14'b00100000111010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00100000111010) && ({row_reg, col_reg}<14'b00100000111101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b00100000111101) && ({row_reg, col_reg}<14'b00100000111111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00100000111111) && ({row_reg, col_reg}<14'b00100001000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00100001000100) && ({row_reg, col_reg}<14'b00100001000110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00100001000110) && ({row_reg, col_reg}<14'b00100010101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b00100010101011) && ({row_reg, col_reg}<14'b00100010101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00100010101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00100010101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00100010110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00100010110001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00100010110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00100010110011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00100010110100) && ({row_reg, col_reg}<14'b00100010110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00100010110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00100010110111) && ({row_reg, col_reg}<14'b00100010111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00100010111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00100010111100) && ({row_reg, col_reg}<14'b00100010111110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00100010111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00100010111111) && ({row_reg, col_reg}<14'b00100011000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00100011000100) && ({row_reg, col_reg}<14'b00100011000110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00100011000110) && ({row_reg, col_reg}<14'b00100100101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00100100101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00100100101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00100100101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00100100101110) && ({row_reg, col_reg}<14'b00100100110000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00100100110000) && ({row_reg, col_reg}<14'b00100100110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00100100110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00100100110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00100100110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00100100110111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00100100111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00100100111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00100100111010) && ({row_reg, col_reg}<14'b00100100111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00100100111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00100100111111) && ({row_reg, col_reg}<14'b00100101000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00100101000010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00100101000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00100101000100)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00100101000101) && ({row_reg, col_reg}<14'b00100110101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00100110101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00100110101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00100110101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00100110101101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00100110101110) && ({row_reg, col_reg}<14'b00100110110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00100110110000) && ({row_reg, col_reg}<14'b00100110110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00100110110011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00100110110100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00100110110101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00100110110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00100110110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b00100110111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b00100110111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00100110111010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00100110111011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00100110111100) && ({row_reg, col_reg}<14'b00100111000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00100111000000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00100111000001) && ({row_reg, col_reg}<14'b00100111000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00100111000100)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00100111000101) && ({row_reg, col_reg}<14'b00101000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b00101000101010) && ({row_reg, col_reg}<14'b00101000101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00101000101101) && ({row_reg, col_reg}<14'b00101000110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00101000110001) && ({row_reg, col_reg}<14'b00101000110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00101000110011) && ({row_reg, col_reg}<14'b00101000110111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00101000110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00101000111000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00101000111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b00101000111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b00101000111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00101000111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00101000111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00101000111110) && ({row_reg, col_reg}<14'b00101001000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00101001000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00101001000001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00101001000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00101001000011) && ({row_reg, col_reg}<14'b00101001000101)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00101001000101) && ({row_reg, col_reg}<14'b00101010101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00101010101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00101010101010) && ({row_reg, col_reg}<14'b00101010101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00101010101101) && ({row_reg, col_reg}<14'b00101010110001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00101010110001) && ({row_reg, col_reg}<14'b00101010110011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00101010110011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00101010110100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00101010110101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00101010110110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00101010110111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00101010111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00101010111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00101010111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00101010111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b00101010111100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00101010111101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00101010111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00101010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00101011000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00101011000001) && ({row_reg, col_reg}<14'b00101011000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00101011000011)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00101011000100) && ({row_reg, col_reg}<14'b00101100101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00101100101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00101100101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00101100101011)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==14'b00101100101100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=14'b00101100101101) && ({row_reg, col_reg}<14'b00101100110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00101100110000) && ({row_reg, col_reg}<14'b00101100110010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00101100110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00101100110011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00101100110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00101100110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b00101100110110) && ({row_reg, col_reg}<14'b00101100111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b00101100111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b00101100111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b00101100111010) && ({row_reg, col_reg}<14'b00101100111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00101100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00101100111101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b00101100111110) && ({row_reg, col_reg}<14'b00101101000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00101101000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00101101000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00101101000010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00101101000011)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00101101000100) && ({row_reg, col_reg}<14'b00101110101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b00101110101000) && ({row_reg, col_reg}<14'b00101110101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00101110101011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b00101110101100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b00101110101101) && ({row_reg, col_reg}<14'b00101110110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00101110110000) && ({row_reg, col_reg}<14'b00101110110010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00101110110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00101110110011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b00101110110100) && ({row_reg, col_reg}<14'b00101110110110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00101110110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00101110110111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00101110111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00101110111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b00101110111010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00101110111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00101110111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00101110111101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00101110111110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00101110111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00101111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00101111000001) && ({row_reg, col_reg}<14'b00101111000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00101111000011)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00101111000100) && ({row_reg, col_reg}<14'b00110000101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b00110000101000) && ({row_reg, col_reg}<14'b00110000101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00110000101010) && ({row_reg, col_reg}<14'b00110000101100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b00110000101100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b00110000101101) && ({row_reg, col_reg}<14'b00110000101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00110000101111) && ({row_reg, col_reg}<14'b00110000110001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00110000110001) && ({row_reg, col_reg}<14'b00110000110011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00110000110011) && ({row_reg, col_reg}<14'b00110000110101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00110000110101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00110000110110) && ({row_reg, col_reg}<14'b00110000111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00110000111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00110000111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00110000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b00110000111011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00110000111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00110000111101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00110000111110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00110000111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00110001000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00110001000001) && ({row_reg, col_reg}<14'b00110001000100)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00110001000100) && ({row_reg, col_reg}<14'b00110010101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00110010101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00110010101001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b00110010101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b00110010101011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==14'b00110010101100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=14'b00110010101101) && ({row_reg, col_reg}<14'b00110010101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00110010101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00110010110000) && ({row_reg, col_reg}<14'b00110010110011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00110010110011) && ({row_reg, col_reg}<14'b00110010110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00110010110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00110010110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00110010110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00110010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00110010111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00110010111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00110010111011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00110010111100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00110010111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00110010111110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00110010111111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00110011000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00110011000001) && ({row_reg, col_reg}<14'b00110011000100)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00110011000100) && ({row_reg, col_reg}<14'b00110100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00110100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00110100101001) && ({row_reg, col_reg}<14'b00110100101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b00110100101011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b00110100101100)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b00110100101101) && ({row_reg, col_reg}<14'b00110100101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00110100101111) && ({row_reg, col_reg}<14'b00110100110001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00110100110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00110100110010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b00110100110011) && ({row_reg, col_reg}<14'b00110100110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00110100110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b00110100110110) && ({row_reg, col_reg}<14'b00110100111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b00110100111000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00110100111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00110100111010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00110100111011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00110100111100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00110100111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00110100111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00110100111111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00110101000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00110101000001) && ({row_reg, col_reg}<14'b00110101000101)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00110101000101) && ({row_reg, col_reg}<14'b00110110101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00110110101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00110110101001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b00110110101010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b00110110101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b00110110101100) && ({row_reg, col_reg}<14'b00110110101110)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==14'b00110110101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00110110101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00110110110000) && ({row_reg, col_reg}<14'b00110110110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00110110110010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00110110110011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00110110110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00110110110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b00110110110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b00110110110111) && ({row_reg, col_reg}<14'b00110110111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b00110110111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b00110110111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b00110110111011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00110110111100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00110110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00110110111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00110110111111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00110111000000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00110111000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00110111000010) && ({row_reg, col_reg}<14'b00110111000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00110111000110)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=14'b00110111000111) && ({row_reg, col_reg}<14'b00111000101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b00111000101001) && ({row_reg, col_reg}<14'b00111000101011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b00111000101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b00111000101100)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b00111000101101) && ({row_reg, col_reg}<14'b00111000101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00111000101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00111000110000) && ({row_reg, col_reg}<14'b00111000110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00111000110010) && ({row_reg, col_reg}<14'b00111000110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00111000110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00111000110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b00111000110110) && ({row_reg, col_reg}<14'b00111000111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b00111000111000) && ({row_reg, col_reg}<14'b00111000111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b00111000111010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00111000111011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00111000111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00111000111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00111000111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00111000111111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00111001000000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00111001000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00111001000010) && ({row_reg, col_reg}<14'b00111001000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00111001000101) && ({row_reg, col_reg}<14'b00111001001000)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=14'b00111001001000) && ({row_reg, col_reg}<14'b00111010101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00111010101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b00111010101010)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==14'b00111010101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b00111010101100)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b00111010101101) && ({row_reg, col_reg}<14'b00111010101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00111010101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00111010110000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00111010110001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00111010110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00111010110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00111010110100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b00111010110101) && ({row_reg, col_reg}<14'b00111010110111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=14'b00111010110111) && ({row_reg, col_reg}<14'b00111010111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b00111010111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b00111010111010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b00111010111011) && ({row_reg, col_reg}<14'b00111010111101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00111010111101) && ({row_reg, col_reg}<14'b00111010111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00111010111111) && ({row_reg, col_reg}<14'b00111011000001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00111011000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00111011000010) && ({row_reg, col_reg}<14'b00111011000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00111011000100) && ({row_reg, col_reg}<14'b00111011001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00111011001000)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00111011001001) && ({row_reg, col_reg}<14'b00111100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00111100101000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b00111100101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b00111100101010)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==14'b00111100101011)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==14'b00111100101100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=14'b00111100101101) && ({row_reg, col_reg}<14'b00111100110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00111100110000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00111100110001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00111100110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b00111100110011) && ({row_reg, col_reg}<14'b00111100110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00111100110101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00111100110110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b00111100110111) && ({row_reg, col_reg}<14'b00111100111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b00111100111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b00111100111010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00111100111011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00111100111100) && ({row_reg, col_reg}<14'b00111100111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00111100111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00111100111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00111101000000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00111101000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00111101000010) && ({row_reg, col_reg}<14'b00111101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00111101000100) && ({row_reg, col_reg}<14'b00111101000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00111101000111) && ({row_reg, col_reg}<14'b00111101001001)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00111101001001) && ({row_reg, col_reg}<14'b00111110101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00111110101000)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b00111110101001) && ({row_reg, col_reg}<14'b00111110101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b00111110101011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b00111110101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00111110101101) && ({row_reg, col_reg}<14'b00111110101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00111110101111) && ({row_reg, col_reg}<14'b00111110110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00111110110001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00111110110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00111110110011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00111110110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00111110110101) && ({row_reg, col_reg}<14'b00111110110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00111110110111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00111110111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b00111110111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b00111110111010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00111110111011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00111110111100) && ({row_reg, col_reg}<14'b00111110111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00111110111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00111110111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00111111000000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00111111000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00111111000010) && ({row_reg, col_reg}<14'b00111111000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00111111000100) && ({row_reg, col_reg}<14'b00111111000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00111111000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00111111001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00111111001001)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00111111001010) && ({row_reg, col_reg}<14'b01000000101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000000101000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==14'b01000000101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000000101010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b01000000101011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b01000000101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01000000101101) && ({row_reg, col_reg}<14'b01000000101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01000000101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01000000110000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01000000110001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01000000110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01000000110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01000000110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b01000000110101) && ({row_reg, col_reg}<14'b01000000110111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01000000110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01000000111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01000000111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01000000111010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01000000111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01000000111100) && ({row_reg, col_reg}<14'b01000000111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01000000111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01000000111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01000001000000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01000001000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01000001000010) && ({row_reg, col_reg}<14'b01000001000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01000001000100) && ({row_reg, col_reg}<14'b01000001000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01000001000111) && ({row_reg, col_reg}<14'b01000001001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01000001001001)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=14'b01000001001010) && ({row_reg, col_reg}<14'b01000010101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000010101001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b01000010101010)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==14'b01000010101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==14'b01000010101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01000010101101) && ({row_reg, col_reg}<14'b01000010101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01000010101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01000010110000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01000010110001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01000010110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01000010110011) && ({row_reg, col_reg}<14'b01000010110111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01000010110111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01000010111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01000010111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01000010111010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01000010111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01000010111100) && ({row_reg, col_reg}<14'b01000010111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01000010111110) && ({row_reg, col_reg}<14'b01000011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01000011000000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01000011000001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01000011000010) && ({row_reg, col_reg}<14'b01000011000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01000011000100) && ({row_reg, col_reg}<14'b01000011000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01000011000111) && ({row_reg, col_reg}<14'b01000011001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01000011001001)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=14'b01000011001010) && ({row_reg, col_reg}<14'b01000100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000100100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b01000100101000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b01000100101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01000100101010)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==14'b01000100101011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==14'b01000100101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01000100101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01000100101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01000100101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01000100110000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b01000100110001) && ({row_reg, col_reg}<14'b01000100110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01000100110011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b01000100110100) && ({row_reg, col_reg}<14'b01000100110111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=14'b01000100110111) && ({row_reg, col_reg}<14'b01000100111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01000100111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01000100111010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01000100111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01000100111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01000100111101) && ({row_reg, col_reg}<14'b01000101000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01000101000000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01000101000001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01000101000010) && ({row_reg, col_reg}<14'b01000101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01000101000100) && ({row_reg, col_reg}<14'b01000101000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01000101000110) && ({row_reg, col_reg}<14'b01000101001011)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b01000101001011) && ({row_reg, col_reg}<14'b01000110100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000110100111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b01000110101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01000110101001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b01000110101010)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==14'b01000110101011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b01000110101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01000110101101) && ({row_reg, col_reg}<14'b01000110101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01000110101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01000110110000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b01000110110001) && ({row_reg, col_reg}<14'b01000110110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01000110110011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b01000110110100) && ({row_reg, col_reg}<14'b01000110110111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01000110110111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01000110111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01000110111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01000110111010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01000110111011) && ({row_reg, col_reg}<14'b01000110111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01000110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01000110111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01000110111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01000111000000) && ({row_reg, col_reg}<14'b01000111000010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01000111000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01000111000011) && ({row_reg, col_reg}<14'b01000111000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01000111000110) && ({row_reg, col_reg}<14'b01000111001011)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b01000111001011) && ({row_reg, col_reg}<14'b01001000100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001000100111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b01001000101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b01001000101001) && ({row_reg, col_reg}<14'b01001000101011)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b01001000101011) && ({row_reg, col_reg}<14'b01001000101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01001000101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01001000101110) && ({row_reg, col_reg}<14'b01001000110000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01001000110000) && ({row_reg, col_reg}<14'b01001000110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01001000110010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01001000110011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b01001000110100) && ({row_reg, col_reg}<14'b01001000110110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01001000110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01001000110111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01001000111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01001000111001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01001000111010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01001000111011) && ({row_reg, col_reg}<14'b01001000111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01001000111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01001000111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01001000111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01001001000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01001001000001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01001001000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01001001000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01001001000100) && ({row_reg, col_reg}<14'b01001001000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01001001000110) && ({row_reg, col_reg}<14'b01001001001011)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b01001001001011) && ({row_reg, col_reg}<14'b01001010100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001010100111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b01001010101000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=14'b01001010101001) && ({row_reg, col_reg}<14'b01001010101011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b01001010101011) && ({row_reg, col_reg}<14'b01001010101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01001010101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01001010101110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01001010101111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01001010110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01001010110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01001010110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01001010110011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b01001010110100) && ({row_reg, col_reg}<14'b01001010110110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01001010110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01001010110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01001010111000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01001010111001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01001010111010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01001010111011) && ({row_reg, col_reg}<14'b01001010111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01001010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01001010111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01001010111111) && ({row_reg, col_reg}<14'b01001011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01001011000001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01001011000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01001011000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01001011000100) && ({row_reg, col_reg}<14'b01001011000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01001011000110) && ({row_reg, col_reg}<14'b01001011001011)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b01001011001011) && ({row_reg, col_reg}<14'b01001100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001100100110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01001100100111)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==14'b01001100101000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b01001100101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01001100101010)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b01001100101011) && ({row_reg, col_reg}<14'b01001100101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01001100101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01001100101110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01001100101111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01001100110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01001100110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01001100110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01001100110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01001100110100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01001100110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01001100110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01001100110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01001100111000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01001100111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01001100111010) && ({row_reg, col_reg}<14'b01001100111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01001100111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01001100111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01001101000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01001101000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01001101000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01001101000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01001101000100) && ({row_reg, col_reg}<14'b01001101000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01001101000110) && ({row_reg, col_reg}<14'b01001101001011)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b01001101001011) && ({row_reg, col_reg}<14'b01001110100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001110100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==14'b01001110100111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b01001110101000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==14'b01001110101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b01001110101010) && ({row_reg, col_reg}<14'b01001110101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01001110101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01001110101101) && ({row_reg, col_reg}<14'b01001110101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01001110101111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b01001110110000) && ({row_reg, col_reg}<14'b01001110110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01001110110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01001110110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01001110110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01001110110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01001110110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01001110111000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01001110111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01001110111010) && ({row_reg, col_reg}<14'b01001110111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01001110111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01001110111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01001110111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01001110111111) && ({row_reg, col_reg}<14'b01001111000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01001111000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01001111000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01001111000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01001111000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01001111000101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01001111000110) && ({row_reg, col_reg}<14'b01001111001100)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b01001111001100) && ({row_reg, col_reg}<14'b01010000100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010000100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b01010000100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010000101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b01010000101001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=14'b01010000101010) && ({row_reg, col_reg}<14'b01010000101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01010000101101) && ({row_reg, col_reg}<14'b01010000101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01010000101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01010000110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01010000110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01010000110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01010000110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01010000110100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01010000110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01010000110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01010000110111) && ({row_reg, col_reg}<14'b01010000111001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01010000111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01010000111010) && ({row_reg, col_reg}<14'b01010000111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01010000111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01010000111101) && ({row_reg, col_reg}<14'b01010000111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01010000111111) && ({row_reg, col_reg}<14'b01010001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01010001000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01010001000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01010001000011) && ({row_reg, col_reg}<14'b01010001000101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01010001000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01010001000110) && ({row_reg, col_reg}<14'b01010001001100)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b01010001001100) && ({row_reg, col_reg}<14'b01010010100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010010100111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b01010010101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01010010101001)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==14'b01010010101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01010010101011) && ({row_reg, col_reg}<14'b01010010101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01010010101101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01010010101110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01010010101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01010010110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01010010110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b01010010110010) && ({row_reg, col_reg}<14'b01010010110100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01010010110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01010010110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01010010110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01010010110111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01010010111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01010010111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01010010111010) && ({row_reg, col_reg}<14'b01010010111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01010010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01010010111101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01010010111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01010010111111) && ({row_reg, col_reg}<14'b01010011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01010011000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01010011000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01010011000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01010011000100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01010011000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01010011000110) && ({row_reg, col_reg}<14'b01010011001100)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b01010011001100) && ({row_reg, col_reg}<14'b01010100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010100100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b01010100100111) && ({row_reg, col_reg}<14'b01010100101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01010100101001)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==14'b01010100101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01010100101011) && ({row_reg, col_reg}<14'b01010100101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01010100101101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01010100101110) && ({row_reg, col_reg}<14'b01010100110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01010100110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01010100110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01010100110010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01010100110011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01010100110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b01010100110101) && ({row_reg, col_reg}<14'b01010100110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01010100110111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01010100111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01010100111001) && ({row_reg, col_reg}<14'b01010100111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01010100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01010100111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01010100111101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01010100111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01010100111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01010101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01010101000001) && ({row_reg, col_reg}<14'b01010101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01010101000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01010101000100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01010101000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01010101000110) && ({row_reg, col_reg}<14'b01010101001100)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b01010101001100) && ({row_reg, col_reg}<14'b01010110100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010110100101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=14'b01010110100110) && ({row_reg, col_reg}<14'b01010110101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b01010110101001) && ({row_reg, col_reg}<14'b01010110101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01010110101011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01010110101100) && ({row_reg, col_reg}<14'b01010110101110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01010110101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01010110101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01010110110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01010110110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b01010110110010) && ({row_reg, col_reg}<14'b01010110110100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01010110110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01010110110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01010110110110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01010110110111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b01010110111000) && ({row_reg, col_reg}<14'b01010110111010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01010110111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01010110111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01010110111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01010110111101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01010110111110) && ({row_reg, col_reg}<14'b01010111000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01010111000000) && ({row_reg, col_reg}<14'b01010111000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01010111000011) && ({row_reg, col_reg}<14'b01010111000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01010111000110) && ({row_reg, col_reg}<14'b01010111001100)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b01010111001100) && ({row_reg, col_reg}<14'b01011000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011000100101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b01011000100110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=14'b01011000100111) && ({row_reg, col_reg}<14'b01011000101001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b01011000101001) && ({row_reg, col_reg}<14'b01011000101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01011000101011) && ({row_reg, col_reg}<14'b01011000101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01011000101101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01011000101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01011000101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01011000110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01011000110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01011000110010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01011000110011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01011000110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01011000110101) && ({row_reg, col_reg}<14'b01011000110111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01011000110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01011000111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01011000111001) && ({row_reg, col_reg}<14'b01011000111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01011000111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01011000111100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01011000111101) && ({row_reg, col_reg}<14'b01011000111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01011000111111) && ({row_reg, col_reg}<14'b01011001000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01011001000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011001000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01011001000100) && ({row_reg, col_reg}<14'b01011001000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01011001000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01011001000111) && ({row_reg, col_reg}<14'b01011001001100)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b01011001001100) && ({row_reg, col_reg}<14'b01011010100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011010100101)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==14'b01011010100110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b01011010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01011010101000)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b01011010101001) && ({row_reg, col_reg}<14'b01011010101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01011010101100) && ({row_reg, col_reg}<14'b01011010101110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01011010101110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01011010101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01011010110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01011010110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01011010110010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01011010110011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01011010110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b01011010110101) && ({row_reg, col_reg}<14'b01011010110111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01011010110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01011010111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01011010111001) && ({row_reg, col_reg}<14'b01011010111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01011010111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01011010111100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01011010111101) && ({row_reg, col_reg}<14'b01011010111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01011010111111) && ({row_reg, col_reg}<14'b01011011000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01011011000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011011000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01011011000100) && ({row_reg, col_reg}<14'b01011011000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01011011000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01011011000111) && ({row_reg, col_reg}<14'b01011011001100)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b01011011001100) && ({row_reg, col_reg}<14'b01011100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011100100100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b01011100100101) && ({row_reg, col_reg}<14'b01011100100111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==14'b01011100100111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b01011100101000)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b01011100101001) && ({row_reg, col_reg}<14'b01011100101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01011100101100) && ({row_reg, col_reg}<14'b01011100101110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01011100101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01011100101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01011100110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b01011100110001) && ({row_reg, col_reg}<14'b01011100110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01011100110011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01011100110100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01011100110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01011100110110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01011100110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01011100111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01011100111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01011100111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01011100111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01011100111100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01011100111101) && ({row_reg, col_reg}<14'b01011100111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01011100111111) && ({row_reg, col_reg}<14'b01011101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01011101000001) && ({row_reg, col_reg}<14'b01011101000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01011101000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01011101000101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01011101000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01011101000111) && ({row_reg, col_reg}<14'b01011101001100)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b01011101001100) && ({row_reg, col_reg}<14'b01011110100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011110100110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b01011110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b01011110101000) && ({row_reg, col_reg}<14'b01011110101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01011110101011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01011110101100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01011110101101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b01011110101110) && ({row_reg, col_reg}<14'b01011110110001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01011110110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01011110110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01011110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011110110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01011110110101) && ({row_reg, col_reg}<14'b01011110110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01011110110111) && ({row_reg, col_reg}<14'b01011110111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01011110111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01011110111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01011110111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01011110111100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01011110111101) && ({row_reg, col_reg}<14'b01011110111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01011110111111) && ({row_reg, col_reg}<14'b01011111000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01011111000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01011111000010) && ({row_reg, col_reg}<14'b01011111000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01011111000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01011111000101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01011111000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01011111000111) && ({row_reg, col_reg}<14'b01011111001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01011111001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01011111001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b01011111001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01011111001111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b01011111010000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b01011111010001)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==14'b01011111010010)) color_data = 12'b010000110001;

		if(({row_reg, col_reg}>=14'b01011111010011) && ({row_reg, col_reg}<14'b01100000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100000100101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=14'b01100000100110) && ({row_reg, col_reg}<14'b01100000101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b01100000101000) && ({row_reg, col_reg}<14'b01100000101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01100000101010) && ({row_reg, col_reg}<14'b01100000101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01100000101100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01100000101101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01100000101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01100000101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01100000110000) && ({row_reg, col_reg}<14'b01100000110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01100000110010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01100000110011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01100000110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100000110101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01100000110110) && ({row_reg, col_reg}<14'b01100000111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01100000111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01100000111001) && ({row_reg, col_reg}<14'b01100000111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01100000111011) && ({row_reg, col_reg}<14'b01100000111101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01100000111101) && ({row_reg, col_reg}<14'b01100000111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100000111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01100001000000) && ({row_reg, col_reg}<14'b01100001000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01100001000010) && ({row_reg, col_reg}<14'b01100001000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100001000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100001000101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01100001000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01100001000111) && ({row_reg, col_reg}<14'b01100001001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100001001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b01100001001100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b01100001001101)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}>=14'b01100001001110) && ({row_reg, col_reg}<14'b01100001010001)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==14'b01100001010001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b01100001010010)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==14'b01100001010011)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==14'b01100001010100)) color_data = 12'b010000110001;

		if(({row_reg, col_reg}>=14'b01100001010101) && ({row_reg, col_reg}<14'b01100010100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100010100100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=14'b01100010100101) && ({row_reg, col_reg}<14'b01100010100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01100010100111)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b01100010101000) && ({row_reg, col_reg}<14'b01100010101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100010101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01100010101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01100010101100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01100010101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01100010101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01100010101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01100010110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01100010110001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01100010110010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01100010110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01100010110100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01100010110101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01100010110110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01100010110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01100010111000) && ({row_reg, col_reg}<14'b01100010111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100010111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01100010111100) && ({row_reg, col_reg}<14'b01100010111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01100010111110) && ({row_reg, col_reg}<14'b01100011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100011000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01100011000001) && ({row_reg, col_reg}<14'b01100011000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100011000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100011000101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01100011000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100011000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100011001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01100011001001) && ({row_reg, col_reg}<14'b01100011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100011001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b01100011001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b01100011001101)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}>=14'b01100011001110) && ({row_reg, col_reg}<14'b01100011010000)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}>=14'b01100011010000) && ({row_reg, col_reg}<14'b01100011010010)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}>=14'b01100011010010) && ({row_reg, col_reg}<14'b01100011010101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b01100011010101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b01100011010110)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}>=14'b01100011010111) && ({row_reg, col_reg}<14'b01100100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100100100011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=14'b01100100100100) && ({row_reg, col_reg}<14'b01100100100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01100100100111)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b01100100101000) && ({row_reg, col_reg}<14'b01100100101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100100101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01100100101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01100100101100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01100100101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b01100100101110) && ({row_reg, col_reg}<14'b01100100110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b01100100110000) && ({row_reg, col_reg}<14'b01100100110010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01100100110010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01100100110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b01100100110100) && ({row_reg, col_reg}<14'b01100100110110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01100100110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01100100110111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01100100111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100100111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100100111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100100111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01100100111100) && ({row_reg, col_reg}<14'b01100100111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01100100111110) && ({row_reg, col_reg}<14'b01100101000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01100101000001) && ({row_reg, col_reg}<14'b01100101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100101000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100101000101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01100101000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100101000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100101001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01100101001001) && ({row_reg, col_reg}<14'b01100101001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100101001011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01100101001100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=14'b01100101001101) && ({row_reg, col_reg}<14'b01100101001111)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==14'b01100101001111)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==14'b01100101010000)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}>=14'b01100101010001) && ({row_reg, col_reg}<14'b01100101010011)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}>=14'b01100101010011) && ({row_reg, col_reg}<14'b01100101010111)) color_data = 12'b010000110001;

		if(({row_reg, col_reg}==14'b01100101010111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=14'b01100110000000) && ({row_reg, col_reg}<14'b01100110100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01100110100011) && ({row_reg, col_reg}<14'b01100110100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b01100110100111) && ({row_reg, col_reg}<14'b01100110101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01100110101001) && ({row_reg, col_reg}<14'b01100110101011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01100110101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01100110101100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01100110101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01100110101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01100110101111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b01100110110000) && ({row_reg, col_reg}<14'b01100110110010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01100110110010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01100110110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01100110110100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01100110110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01100110110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01100110110111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01100110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100110111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100110111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100110111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01100110111100) && ({row_reg, col_reg}<14'b01100110111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01100110111110) && ({row_reg, col_reg}<14'b01100111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100111000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100111000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100111000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100111000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100111000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100111000101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01100111000110) && ({row_reg, col_reg}<14'b01100111001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100111001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01100111001001) && ({row_reg, col_reg}<14'b01100111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100111001011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b01100111001100)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}>=14'b01100111001101) && ({row_reg, col_reg}<14'b01100111001111)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==14'b01100111001111)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==14'b01100111010000)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==14'b01100111010001)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==14'b01100111010010)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==14'b01100111010011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b01100111010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b01100111010101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b01100111010110)) color_data = 12'b010000100001;

		if(({row_reg, col_reg}==14'b01100111010111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=14'b01101000000000) && ({row_reg, col_reg}<14'b01101000100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101000100011)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==14'b01101000100100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=14'b01101000100101) && ({row_reg, col_reg}<14'b01101000100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b01101000100111) && ({row_reg, col_reg}<14'b01101000101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101000101001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01101000101010) && ({row_reg, col_reg}<14'b01101000101100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01101000101100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01101000101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01101000101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01101000101111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b01101000110000) && ({row_reg, col_reg}<14'b01101000110010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01101000110010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01101000110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b01101000110100) && ({row_reg, col_reg}<14'b01101000110110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01101000110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01101000110111) && ({row_reg, col_reg}<14'b01101000111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101000111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101000111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101000111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01101000111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101000111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101000111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101000111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01101001000000) && ({row_reg, col_reg}<14'b01101001000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101001000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101001000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01101001000100) && ({row_reg, col_reg}<14'b01101001000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01101001000110) && ({row_reg, col_reg}<14'b01101001001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101001001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101001001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==14'b01101001001011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b01101001001100)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==14'b01101001001101)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}>=14'b01101001001110) && ({row_reg, col_reg}<14'b01101001010001)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==14'b01101001010001)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==14'b01101001010010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b01101001010011)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==14'b01101001010100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01101001010101)) color_data = 12'b010000100001;

		if(({row_reg, col_reg}>=14'b01101001010110) && ({row_reg, col_reg}<14'b01101010000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b01101010000000) && ({row_reg, col_reg}<14'b01101010100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101010100010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b01101010100011)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==14'b01101010100100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b01101010100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01101010100110)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b01101010100111) && ({row_reg, col_reg}<14'b01101010101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101010101001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01101010101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01101010101011) && ({row_reg, col_reg}<14'b01101010101101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01101010101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01101010101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01101010101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01101010110000) && ({row_reg, col_reg}<14'b01101010110010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01101010110010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01101010110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01101010110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01101010110101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01101010110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01101010110111) && ({row_reg, col_reg}<14'b01101010111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101010111010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01101010111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01101010111100) && ({row_reg, col_reg}<14'b01101010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01101011000000) && ({row_reg, col_reg}<14'b01101011000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101011000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101011000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01101011000100) && ({row_reg, col_reg}<14'b01101011000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01101011000110) && ({row_reg, col_reg}<14'b01101011001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01101011001000) && ({row_reg, col_reg}<14'b01101011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101011001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b01101011001011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=14'b01101011001100) && ({row_reg, col_reg}<14'b01101011001110)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}>=14'b01101011001110) && ({row_reg, col_reg}<14'b01101011010001)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==14'b01101011010001)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==14'b01101011010010)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}>=14'b01101011010011) && ({row_reg, col_reg}<14'b01101011010111)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}==14'b01101011010111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=14'b01101100000000) && ({row_reg, col_reg}<14'b01101100100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101100100010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b01101100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101100100100)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==14'b01101100100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b01101100100110) && ({row_reg, col_reg}<14'b01101100101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01101100101000) && ({row_reg, col_reg}<14'b01101100101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01101100101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01101100101011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01101100101100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b01101100101101) && ({row_reg, col_reg}<14'b01101100101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01101100101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101100110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101100110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101100110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01101100110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01101100110100) && ({row_reg, col_reg}<14'b01101100110110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01101100110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01101100110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101100111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101100111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101100111010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01101100111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01101100111100) && ({row_reg, col_reg}<14'b01101100111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101101000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101101000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01101101000010) && ({row_reg, col_reg}<14'b01101101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101101000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01101101000101) && ({row_reg, col_reg}<14'b01101101001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101101001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101101001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b01101101001011)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}>=14'b01101101001100) && ({row_reg, col_reg}<14'b01101101010000)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==14'b01101101010000)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==14'b01101101010001)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==14'b01101101010010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=14'b01101101010011) && ({row_reg, col_reg}<14'b01101101010101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b01101101010101) && ({row_reg, col_reg}<14'b01101101010111)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}>=14'b01101101010111) && ({row_reg, col_reg}<14'b01101110100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101110100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b01101110100011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==14'b01101110100100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b01101110100101)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b01101110100110) && ({row_reg, col_reg}<14'b01101110101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101110101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01101110101001) && ({row_reg, col_reg}<14'b01101110101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01101110101011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01101110101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01101110101101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01101110101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01101110101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01101110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101110110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101110110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101110110011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01101110110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01101110110101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01101110110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01101110110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101110111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101110111010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01101110111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101110111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101110111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01101110111110) && ({row_reg, col_reg}<14'b01101111000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101111000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101111000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101111000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101111000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01101111000101) && ({row_reg, col_reg}<14'b01101111001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01101111001000) && ({row_reg, col_reg}<14'b01101111001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101111001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b01101111001011)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}>=14'b01101111001100) && ({row_reg, col_reg}<14'b01101111010000)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==14'b01101111010000)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==14'b01101111010001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b01101111010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b01101111010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b01101111010100) && ({row_reg, col_reg}<14'b01101111010110)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}>=14'b01101111010110) && ({row_reg, col_reg}<14'b01110000100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110000100010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==14'b01110000100011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b01110000100100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01110000100101)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b01110000100110) && ({row_reg, col_reg}<14'b01110000101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110000101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01110000101001) && ({row_reg, col_reg}<14'b01110000101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01110000101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01110000101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01110000101101) && ({row_reg, col_reg}<14'b01110000110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01110000110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01110000110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01110000110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110000110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110000110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01110000110101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01110000110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01110000110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110000111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110000111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110000111010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01110000111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110000111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110000111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110000111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01110000111111) && ({row_reg, col_reg}<14'b01110001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110001000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110001000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110001000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110001000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01110001000101) && ({row_reg, col_reg}<14'b01110001001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110001001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01110001001011)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}>=14'b01110001001100) && ({row_reg, col_reg}<14'b01110001010000)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==14'b01110001010000)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==14'b01110001010001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b01110001010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b01110001010011)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}>=14'b01110001010100) && ({row_reg, col_reg}<14'b01110010100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110010100001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==14'b01110010100010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b01110010100011) && ({row_reg, col_reg}<14'b01110010100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b01110010100101) && ({row_reg, col_reg}<14'b01110010101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110010101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01110010101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01110010101010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01110010101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01110010101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01110010101101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01110010101110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01110010101111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01110010110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01110010110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01110010110010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01110010110011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01110010110100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01110010110101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01110010110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01110010110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110010111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01110010111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110010111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110010111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110010111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01110010111111) && ({row_reg, col_reg}<14'b01110011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110011000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110011000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110011000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110011000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01110011000101) && ({row_reg, col_reg}<14'b01110011001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110011001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110011001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110011001010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b01110011001011)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}>=14'b01110011001100) && ({row_reg, col_reg}<14'b01110011001111)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==14'b01110011001111)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==14'b01110011010000)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==14'b01110011010001)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==14'b01110011010010)) color_data = 12'b010000100001;

		if(({row_reg, col_reg}>=14'b01110011010011) && ({row_reg, col_reg}<14'b01110100100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110100100001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b01110100100010) && ({row_reg, col_reg}<14'b01110100100101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01110100100101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01110100100110) && ({row_reg, col_reg}<14'b01110100101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110100101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01110100101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01110100101010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01110100101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01110100101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01110100101101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01110100101110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01110100101111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01110100110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01110100110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01110100110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01110100110011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01110100110100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01110100110101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01110100110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110100110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110100111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110100111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01110100111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110100111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01110100111101) && ({row_reg, col_reg}<14'b01110101000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110101000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01110101000001) && ({row_reg, col_reg}<14'b01110101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01110101000011) && ({row_reg, col_reg}<14'b01110101000101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01110101000101) && ({row_reg, col_reg}<14'b01110101001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110101001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110101001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110101001010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b01110101001011)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}>=14'b01110101001100) && ({row_reg, col_reg}<14'b01110101001110)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}>=14'b01110101001110) && ({row_reg, col_reg}<14'b01110101010000)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==14'b01110101010000)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==14'b01110101010001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b01110101010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01110101010011)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}>=14'b01110101010100) && ({row_reg, col_reg}<14'b01110110100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01110110100001) && ({row_reg, col_reg}<14'b01110110100100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01110110100100)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b01110110100101) && ({row_reg, col_reg}<14'b01110110101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110110101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01110110101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01110110101010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01110110101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01110110101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01110110101101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01110110101110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01110110101111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01110110110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01110110110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01110110110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01110110110011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01110110110100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01110110110101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01110110110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110110110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110110111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01110110111010) && ({row_reg, col_reg}<14'b01110110111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01110110111101) && ({row_reg, col_reg}<14'b01110111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110111000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01110111000001) && ({row_reg, col_reg}<14'b01110111000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01110111000101) && ({row_reg, col_reg}<14'b01110111001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110111001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b01110111001010)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}>=14'b01110111001011) && ({row_reg, col_reg}<14'b01110111001111)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==14'b01110111001111)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==14'b01110111010000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b01110111010001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b01110111010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01110111010011)) color_data = 12'b010000110001;

		if(({row_reg, col_reg}>=14'b01110111010100) && ({row_reg, col_reg}<14'b01111000100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01111000100001) && ({row_reg, col_reg}<14'b01111000100100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01111000100100)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b01111000100101) && ({row_reg, col_reg}<14'b01111000101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111000101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01111000101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01111000101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01111000101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01111000101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01111000101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b01111000101110) && ({row_reg, col_reg}<14'b01111000110000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01111000110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01111000110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01111000110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01111000110011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01111000110100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01111000110101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01111000110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111000110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111000111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111000111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01111000111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111000111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01111000111100) && ({row_reg, col_reg}<14'b01111001000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111001000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01111001000001) && ({row_reg, col_reg}<14'b01111001000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111001000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01111001000110) && ({row_reg, col_reg}<14'b01111001001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111001001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01111001001010)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==14'b01111001001011)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}>=14'b01111001001100) && ({row_reg, col_reg}<14'b01111001001110)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==14'b01111001001110)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==14'b01111001001111)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==14'b01111001010000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b01111001010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01111001010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b01111001010011)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==14'b01111001010100)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}>=14'b01111001010101) && ({row_reg, col_reg}<14'b01111010100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111010100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b01111010100001) && ({row_reg, col_reg}<14'b01111010100011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b01111010100011)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b01111010100100) && ({row_reg, col_reg}<14'b01111010100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111010100111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01111010101000) && ({row_reg, col_reg}<14'b01111010101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01111010101010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01111010101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01111010101100) && ({row_reg, col_reg}<14'b01111010101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b01111010101110) && ({row_reg, col_reg}<14'b01111010110001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01111010110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01111010110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01111010110011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01111010110100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01111010110101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01111010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01111010110111) && ({row_reg, col_reg}<14'b01111010111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111010111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111010111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01111010111100) && ({row_reg, col_reg}<14'b01111011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111011000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01111011000001) && ({row_reg, col_reg}<14'b01111011000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111011000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01111011000111) && ({row_reg, col_reg}<14'b01111011001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111011001001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b01111011001010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=14'b01111011001011) && ({row_reg, col_reg}<14'b01111011001101)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}>=14'b01111011001101) && ({row_reg, col_reg}<14'b01111011001111)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==14'b01111011001111)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==14'b01111011010000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b01111011010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01111011010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b01111011010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b01111011010100)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}>=14'b01111011010101) && ({row_reg, col_reg}<14'b01111100100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111100100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b01111100100001) && ({row_reg, col_reg}<14'b01111100100011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b01111100100011)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b01111100100100) && ({row_reg, col_reg}<14'b01111100100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111100100111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01111100101000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01111100101001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01111100101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01111100101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01111100101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01111100101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01111100101110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01111100101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b01111100110000) && ({row_reg, col_reg}<14'b01111100110010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01111100110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01111100110011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01111100110100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01111100110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111100110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111100111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01111100111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01111100111010) && ({row_reg, col_reg}<14'b01111100111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01111100111111) && ({row_reg, col_reg}<14'b01111101000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01111101000001) && ({row_reg, col_reg}<14'b01111101001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111101001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b01111101001001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=14'b01111101001010) && ({row_reg, col_reg}<14'b01111101001100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=14'b01111101001100) && ({row_reg, col_reg}<14'b01111101010000)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}>=14'b01111101010000) && ({row_reg, col_reg}<14'b01111101010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b01111101010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b01111101010011) && ({row_reg, col_reg}<14'b01111101010101)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}>=14'b01111101010101) && ({row_reg, col_reg}<14'b01111110100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01111110100000) && ({row_reg, col_reg}<14'b01111110100010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==14'b01111110100010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b01111110100011)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b01111110100100) && ({row_reg, col_reg}<14'b01111110100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111110100111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01111110101000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01111110101001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01111110101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b01111110101011) && ({row_reg, col_reg}<14'b01111110101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01111110101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01111110101110) && ({row_reg, col_reg}<14'b01111110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111110110001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01111110110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01111110110011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01111110110100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01111110110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111110110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111110110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111110111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01111110111001) && ({row_reg, col_reg}<14'b01111110111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01111110111011) && ({row_reg, col_reg}<14'b01111110111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111110111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01111111000000) && ({row_reg, col_reg}<14'b01111111000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01111111000101) && ({row_reg, col_reg}<14'b01111111000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b01111111001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b01111111001001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=14'b01111111001010) && ({row_reg, col_reg}<14'b01111111001101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=14'b01111111001101) && ({row_reg, col_reg}<14'b01111111001111)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==14'b01111111001111)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==14'b01111111010000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b01111111010001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b01111111010010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b01111111010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b01111111010100)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=14'b01111111010101) && ({row_reg, col_reg}<14'b10000000011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000000011111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==14'b10000000100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10000000100001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=14'b10000000100010) && ({row_reg, col_reg}<14'b10000000100100)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b10000000100100) && ({row_reg, col_reg}<14'b10000000100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10000000100111) && ({row_reg, col_reg}<14'b10000000101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10000000101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10000000101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10000000101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10000000101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10000000101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10000000101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10000000101111) && ({row_reg, col_reg}<14'b10000000110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000000110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10000000110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10000000110011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10000000110100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10000000110101) && ({row_reg, col_reg}<14'b10000000111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10000000111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10000000111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000000111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10000000111011) && ({row_reg, col_reg}<14'b10000000111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000000111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10000001000000) && ({row_reg, col_reg}<14'b10000001000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000001000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000001000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10000001000110) && ({row_reg, col_reg}<14'b10000001001000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10000001001000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10000001001001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b10000001001010)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}>=14'b10000001001011) && ({row_reg, col_reg}<14'b10000001010000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b10000001010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b10000001010001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=14'b10000001010010) && ({row_reg, col_reg}<14'b10000001010100)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=14'b10000001010100) && ({row_reg, col_reg}<14'b10000010011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000010011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b10000010100000) && ({row_reg, col_reg}<14'b10000010100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10000010100010)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b10000010100011) && ({row_reg, col_reg}<14'b10000010100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10000010100111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10000010101000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10000010101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10000010101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b10000010101011) && ({row_reg, col_reg}<14'b10000010101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10000010101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10000010101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10000010101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b10000010110000) && ({row_reg, col_reg}<14'b10000010110010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10000010110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10000010110011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10000010110100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10000010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000010110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10000010110111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10000010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10000010111001) && ({row_reg, col_reg}<14'b10000010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000010111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10000011000000) && ({row_reg, col_reg}<14'b10000011000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000011000101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==14'b10000011000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10000011000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10000011001000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=14'b10000011001001) && ({row_reg, col_reg}<14'b10000011001011)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}>=14'b10000011001011) && ({row_reg, col_reg}<14'b10000011001110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b10000011001110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b10000011001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10000011010000)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==14'b10000011010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b10000011010010) && ({row_reg, col_reg}<14'b10000011010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==14'b10000011010100)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=14'b10000011010101) && ({row_reg, col_reg}<14'b10000100011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000100011110)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=14'b10000100011111) && ({row_reg, col_reg}<14'b10000100100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10000100100010)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b10000100100011) && ({row_reg, col_reg}<14'b10000100100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10000100100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10000100100111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10000100101000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10000100101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10000100101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10000100101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10000100101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b10000100101101) && ({row_reg, col_reg}<14'b10000100101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10000100101111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10000100110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10000100110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10000100110010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10000100110011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10000100110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10000100110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000100110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10000100110111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10000100111000) && ({row_reg, col_reg}<14'b10000100111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10000100111010) && ({row_reg, col_reg}<14'b10000100111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10000100111110) && ({row_reg, col_reg}<14'b10000101000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10000101000000) && ({row_reg, col_reg}<14'b10000101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000101000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000101000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10000101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10000101000111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=14'b10000101001000) && ({row_reg, col_reg}<14'b10000101001100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b10000101001100)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}>=14'b10000101001101) && ({row_reg, col_reg}<14'b10000101001111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=14'b10000101001111) && ({row_reg, col_reg}<14'b10000101010001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b10000101010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=14'b10000101010010) && ({row_reg, col_reg}<14'b10000101010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==14'b10000101010100)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}>=14'b10000101010101) && ({row_reg, col_reg}<14'b10000110011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000110011110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=14'b10000110011111) && ({row_reg, col_reg}<14'b10000110100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10000110100010)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b10000110100011) && ({row_reg, col_reg}<14'b10000110100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10000110100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10000110100111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10000110101000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10000110101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10000110101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10000110101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10000110101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b10000110101101) && ({row_reg, col_reg}<14'b10000110101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b10000110101111) && ({row_reg, col_reg}<14'b10000110110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10000110110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10000110110010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10000110110011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10000110110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10000110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000110110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10000110110111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10000110111000) && ({row_reg, col_reg}<14'b10000110111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10000110111010) && ({row_reg, col_reg}<14'b10000110111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10000110111110) && ({row_reg, col_reg}<14'b10000111000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10000111000000) && ({row_reg, col_reg}<14'b10000111000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000111000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10000111000110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b10000111000111)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}>=14'b10000111001000) && ({row_reg, col_reg}<14'b10000111001101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=14'b10000111001101) && ({row_reg, col_reg}<14'b10000111001111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=14'b10000111001111) && ({row_reg, col_reg}<14'b10000111010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10000111010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10000111010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000111010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=14'b10000111010100) && ({row_reg, col_reg}<14'b10000111010110)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}>=14'b10000111010110) && ({row_reg, col_reg}<14'b10001000011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10001000011110) && ({row_reg, col_reg}<14'b10001000100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b10001000100010) && ({row_reg, col_reg}<14'b10001000100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001000100101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10001000100110) && ({row_reg, col_reg}<14'b10001000101000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10001000101000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10001000101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10001000101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10001000101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10001000101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b10001000101101) && ({row_reg, col_reg}<14'b10001000110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10001000110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10001000110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10001000110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10001000110011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10001000110100) && ({row_reg, col_reg}<14'b10001000111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10001000111010) && ({row_reg, col_reg}<14'b10001000111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001000111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10001000111111) && ({row_reg, col_reg}<14'b10001001000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001001000100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==14'b10001001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10001001000110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b10001001000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b10001001001000)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}>=14'b10001001001001) && ({row_reg, col_reg}<14'b10001001001011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b10001001001011)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==14'b10001001001100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=14'b10001001001101) && ({row_reg, col_reg}<14'b10001001001111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=14'b10001001001111) && ({row_reg, col_reg}<14'b10001001010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10001001010001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=14'b10001001010010) && ({row_reg, col_reg}<14'b10001001010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001001010100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10001001010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10001001010110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=14'b10001001010111) && ({row_reg, col_reg}<14'b10001010011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10001010011110) && ({row_reg, col_reg}<14'b10001010100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10001010100001)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b10001010100010) && ({row_reg, col_reg}<14'b10001010100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001010100101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10001010100110) && ({row_reg, col_reg}<14'b10001010101000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10001010101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10001010101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b10001010101010) && ({row_reg, col_reg}<14'b10001010101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10001010101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b10001010101101) && ({row_reg, col_reg}<14'b10001010101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10001010101111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10001010110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10001010110001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10001010110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10001010110011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10001010110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001010110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001010110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10001010110111) && ({row_reg, col_reg}<14'b10001010111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10001010111010) && ({row_reg, col_reg}<14'b10001010111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001010111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10001010111111) && ({row_reg, col_reg}<14'b10001011000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001011000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10001011000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10001011000110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b10001011000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=14'b10001011001000) && ({row_reg, col_reg}<14'b10001011001100)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==14'b10001011001100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=14'b10001011001101) && ({row_reg, col_reg}<14'b10001011001111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b10001011001111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b10001011010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10001011010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b10001011010010) && ({row_reg, col_reg}<14'b10001011010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001011010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==14'b10001011010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10001011010110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=14'b10001011010111) && ({row_reg, col_reg}<14'b10001100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001100011101)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==14'b10001100011110)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==14'b10001100011111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=14'b10001100100000) && ({row_reg, col_reg}<14'b10001100100010)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b10001100100010) && ({row_reg, col_reg}<14'b10001100100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001100100101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10001100100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10001100100111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10001100101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b10001100101001) && ({row_reg, col_reg}<14'b10001100101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10001100101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10001100101101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10001100101110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10001100101111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10001100110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10001100110001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10001100110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10001100110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001100110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001100110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001100110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10001100110111) && ({row_reg, col_reg}<14'b10001100111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10001100111010) && ({row_reg, col_reg}<14'b10001100111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001100111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10001100111111) && ({row_reg, col_reg}<14'b10001101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001101000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10001101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10001101000110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b10001101000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=14'b10001101001000) && ({row_reg, col_reg}<14'b10001101001011)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==14'b10001101001011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b10001101001100)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}>=14'b10001101001101) && ({row_reg, col_reg}<14'b10001101010000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b10001101010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10001101010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=14'b10001101010010) && ({row_reg, col_reg}<14'b10001101010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001101010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10001101010110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=14'b10001101010111) && ({row_reg, col_reg}<14'b10001110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001110011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10001110011110)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==14'b10001110011111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b10001110100000)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b10001110100001) && ({row_reg, col_reg}<14'b10001110100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001110100101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10001110100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10001110100111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10001110101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10001110101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10001110101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10001110101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10001110101100) && ({row_reg, col_reg}<14'b10001110101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001110101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10001110101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10001110110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10001110110001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10001110110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10001110110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001110110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10001110110101) && ({row_reg, col_reg}<14'b10001110110111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10001110110111) && ({row_reg, col_reg}<14'b10001110111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10001110111010) && ({row_reg, col_reg}<14'b10001110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10001110111101) && ({row_reg, col_reg}<14'b10001110111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10001110111111) && ({row_reg, col_reg}<14'b10001111000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10001111000100) && ({row_reg, col_reg}<14'b10001111000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10001111000110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b10001111000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=14'b10001111001000) && ({row_reg, col_reg}<14'b10001111001011)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}>=14'b10001111001011) && ({row_reg, col_reg}<14'b10001111001101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=14'b10001111001101) && ({row_reg, col_reg}<14'b10001111010000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b10001111010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10001111010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=14'b10001111010010) && ({row_reg, col_reg}<14'b10001111010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10001111010101) && ({row_reg, col_reg}<14'b10001111010111)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=14'b10001111010111) && ({row_reg, col_reg}<14'b10010000011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010000011101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==14'b10010000011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010000011111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b10010000100000)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==14'b10010000100001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10010000100010) && ({row_reg, col_reg}<14'b10010000100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10010000100101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10010000100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10010000100111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10010000101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10010000101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10010000101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10010000101011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10010000101100) && ({row_reg, col_reg}<14'b10010000101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010000101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10010000101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10010000110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10010000110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10010000110010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10010000110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10010000110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10010000110101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10010000110110) && ({row_reg, col_reg}<14'b10010000111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10010000111010) && ({row_reg, col_reg}<14'b10010000111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10010000111101) && ({row_reg, col_reg}<14'b10010000111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10010000111111) && ({row_reg, col_reg}<14'b10010001000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10010001000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==14'b10010001000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b10010001000101) && ({row_reg, col_reg}<14'b10010001000111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b10010001000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=14'b10010001001000) && ({row_reg, col_reg}<14'b10010001001011)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}>=14'b10010001001011) && ({row_reg, col_reg}<14'b10010001001101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=14'b10010001001101) && ({row_reg, col_reg}<14'b10010001010000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b10010001010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10010001010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=14'b10010001010010) && ({row_reg, col_reg}<14'b10010001010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010001010101)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b10010001010110) && ({row_reg, col_reg}<14'b10010010011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010010011101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==14'b10010010011110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b10010010011111)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==14'b10010010100000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=14'b10010010100001) && ({row_reg, col_reg}<14'b10010010100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10010010100011) && ({row_reg, col_reg}<14'b10010010100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10010010100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10010010100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10010010100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10010010101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10010010101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10010010101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10010010101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10010010101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10010010101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10010010101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010010101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10010010110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10010010110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10010010110010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10010010110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10010010110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10010010110101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10010010110110) && ({row_reg, col_reg}<14'b10010010111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10010010111001) && ({row_reg, col_reg}<14'b10010010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10010010111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10010010111110) && ({row_reg, col_reg}<14'b10010011000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10010011000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10010011000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10010011000101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b10010011000110)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==14'b10010011000111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=14'b10010011001000) && ({row_reg, col_reg}<14'b10010011001011)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==14'b10010011001011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b10010011001100)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}>=14'b10010011001101) && ({row_reg, col_reg}<14'b10010011001111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b10010011001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10010011010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10010011010001)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b10010011010010) && ({row_reg, col_reg}<14'b10010100011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010100011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b10010100011101) && ({row_reg, col_reg}<14'b10010100011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10010100011111)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b10010100100000) && ({row_reg, col_reg}<14'b10010100100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10010100100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10010100100011) && ({row_reg, col_reg}<14'b10010100100101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10010100100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10010100100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10010100100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10010100101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10010100101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10010100101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10010100101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10010100101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10010100101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10010100101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10010100101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10010100110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10010100110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10010100110010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10010100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10010100110100) && ({row_reg, col_reg}<14'b10010100110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10010100110110) && ({row_reg, col_reg}<14'b10010100111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10010100111001) && ({row_reg, col_reg}<14'b10010100111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10010100111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10010100111110) && ({row_reg, col_reg}<14'b10010101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10010101000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10010101000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10010101000101)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b10010101000110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b10010101000111)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}>=14'b10010101001000) && ({row_reg, col_reg}<14'b10010101001100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=14'b10010101001100) && ({row_reg, col_reg}<14'b10010101001110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b10010101001110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b10010101001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10010101010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10010101010001)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b10010101010010) && ({row_reg, col_reg}<14'b10010110011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010110011100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=14'b10010110011101) && ({row_reg, col_reg}<14'b10010110011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10010110011111)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b10010110100000) && ({row_reg, col_reg}<14'b10010110100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10010110100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10010110100011) && ({row_reg, col_reg}<14'b10010110100101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10010110100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10010110100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10010110100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10010110101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10010110101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b10010110101010) && ({row_reg, col_reg}<14'b10010110101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10010110101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10010110101101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b10010110101110) && ({row_reg, col_reg}<14'b10010110110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10010110110000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10010110110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10010110110010) && ({row_reg, col_reg}<14'b10010110110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10010110110100) && ({row_reg, col_reg}<14'b10010110110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10010110110110) && ({row_reg, col_reg}<14'b10010110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10010110111000) && ({row_reg, col_reg}<14'b10010110111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10010110111100) && ({row_reg, col_reg}<14'b10010110111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10010110111110) && ({row_reg, col_reg}<14'b10010111000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10010111000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10010111000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10010111000101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=14'b10010111000110) && ({row_reg, col_reg}<14'b10010111001000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=14'b10010111001000) && ({row_reg, col_reg}<14'b10010111001010)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}>=14'b10010111001010) && ({row_reg, col_reg}<14'b10010111001100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=14'b10010111001100) && ({row_reg, col_reg}<14'b10010111001110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=14'b10010111001110) && ({row_reg, col_reg}<14'b10010111010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10010111010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10010111010001)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b10010111010010) && ({row_reg, col_reg}<14'b10011000011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011000011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10011000011100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=14'b10011000011101) && ({row_reg, col_reg}<14'b10011000011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10011000011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10011000100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10011000100001) && ({row_reg, col_reg}<14'b10011000100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10011000100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10011000100100) && ({row_reg, col_reg}<14'b10011000100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10011000100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10011000100111) && ({row_reg, col_reg}<14'b10011000101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b10011000101001) && ({row_reg, col_reg}<14'b10011000101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b10011000101011) && ({row_reg, col_reg}<14'b10011000101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10011000101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10011000101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10011000110000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10011000110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10011000110010) && ({row_reg, col_reg}<14'b10011000110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10011000110100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10011000110101) && ({row_reg, col_reg}<14'b10011000111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10011000111000) && ({row_reg, col_reg}<14'b10011000111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10011000111100) && ({row_reg, col_reg}<14'b10011000111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10011000111110) && ({row_reg, col_reg}<14'b10011001000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10011001000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b10011001000011) && ({row_reg, col_reg}<14'b10011001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10011001000101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=14'b10011001000110) && ({row_reg, col_reg}<14'b10011001001001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b10011001001001)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==14'b10011001001010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b10011001001011)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==14'b10011001001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b10011001001101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=14'b10011001001110) && ({row_reg, col_reg}<14'b10011001010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10011001010000)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b10011001010001) && ({row_reg, col_reg}<14'b10011010011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10011010011011) && ({row_reg, col_reg}<14'b10011010011101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b10011010011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10011010011110)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b10011010011111) && ({row_reg, col_reg}<14'b10011010100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10011010100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10011010100100) && ({row_reg, col_reg}<14'b10011010100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10011010100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10011010100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b10011010101000) && ({row_reg, col_reg}<14'b10011010101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b10011010101011) && ({row_reg, col_reg}<14'b10011010101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10011010101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10011010101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10011010110000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10011010110001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10011010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10011010110011) && ({row_reg, col_reg}<14'b10011010110101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10011010110101) && ({row_reg, col_reg}<14'b10011010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10011010111000) && ({row_reg, col_reg}<14'b10011010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10011010111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10011010111101) && ({row_reg, col_reg}<14'b10011011000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10011011000010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=14'b10011011000011) && ({row_reg, col_reg}<14'b10011011000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b10011011000101) && ({row_reg, col_reg}<14'b10011011001010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=14'b10011011001010) && ({row_reg, col_reg}<14'b10011011001100)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==14'b10011011001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=14'b10011011001101) && ({row_reg, col_reg}<14'b10011011001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10011011001111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10011011010000)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b10011011010001) && ({row_reg, col_reg}<14'b10011100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10011100011010) && ({row_reg, col_reg}<14'b10011100011100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=14'b10011100011100) && ({row_reg, col_reg}<14'b10011100011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10011100011110)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b10011100011111) && ({row_reg, col_reg}<14'b10011100100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10011100100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10011100100100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10011100100101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10011100100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10011100100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10011100101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b10011100101001) && ({row_reg, col_reg}<14'b10011100101011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10011100101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10011100101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b10011100101101) && ({row_reg, col_reg}<14'b10011100101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10011100101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10011100110000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10011100110001) && ({row_reg, col_reg}<14'b10011100110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10011100110011) && ({row_reg, col_reg}<14'b10011100110101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10011100110101) && ({row_reg, col_reg}<14'b10011100111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10011100111000) && ({row_reg, col_reg}<14'b10011100111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10011100111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10011100111101) && ({row_reg, col_reg}<14'b10011101000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10011101000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b10011101000011) && ({row_reg, col_reg}<14'b10011101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b10011101000101) && ({row_reg, col_reg}<14'b10011101001010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b10011101001010)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==14'b10011101001011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=14'b10011101001100) && ({row_reg, col_reg}<14'b10011101001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10011101001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10011101010000)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b10011101010001) && ({row_reg, col_reg}<14'b10011110011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011110011010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b10011110011011)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}>=14'b10011110011100) && ({row_reg, col_reg}<14'b10011110011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b10011110011110) && ({row_reg, col_reg}<14'b10011110100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10011110100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10011110100011) && ({row_reg, col_reg}<14'b10011110100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10011110100101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10011110100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10011110100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10011110101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b10011110101001) && ({row_reg, col_reg}<14'b10011110101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10011110101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10011110101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10011110101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10011110101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10011110101111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10011110110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10011110110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10011110110010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10011110110011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10011110110100) && ({row_reg, col_reg}<14'b10011110110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10011110110111) && ({row_reg, col_reg}<14'b10011110111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10011110111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10011110111101) && ({row_reg, col_reg}<14'b10011111000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10011111000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=14'b10011111000011) && ({row_reg, col_reg}<14'b10011111000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10011111000101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b10011111000110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b10011111000111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=14'b10011111001000) && ({row_reg, col_reg}<14'b10011111001011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b10011111001011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=14'b10011111001100) && ({row_reg, col_reg}<14'b10011111001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10011111001111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10011111010000)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b10011111010001) && ({row_reg, col_reg}<14'b10100000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10100000011001) && ({row_reg, col_reg}<14'b10100000011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10100000011011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==14'b10100000011100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b10100000011101)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b10100000011110) && ({row_reg, col_reg}<14'b10100000100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10100000100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10100000100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10100000100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10100000100101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b10100000100110) && ({row_reg, col_reg}<14'b10100000101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10100000101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10100000101001) && ({row_reg, col_reg}<14'b10100000101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100000101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10100000101100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10100000101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10100000101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10100000101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10100000110000) && ({row_reg, col_reg}<14'b10100000110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10100000110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10100000110011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10100000110100) && ({row_reg, col_reg}<14'b10100000110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10100000110111) && ({row_reg, col_reg}<14'b10100000111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10100000111011) && ({row_reg, col_reg}<14'b10100000111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10100000111101) && ({row_reg, col_reg}<14'b10100001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10100001000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10100001000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=14'b10100001000011) && ({row_reg, col_reg}<14'b10100001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10100001000110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=14'b10100001000111) && ({row_reg, col_reg}<14'b10100001001011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=14'b10100001001011) && ({row_reg, col_reg}<14'b10100001001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10100001001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10100001001111)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=14'b10100001010000) && ({row_reg, col_reg}<14'b10100010011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10100010011001) && ({row_reg, col_reg}<14'b10100010011100)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==14'b10100010011100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=14'b10100010011101) && ({row_reg, col_reg}<14'b10100010100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10100010100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10100010100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10100010100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10100010100101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10100010100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10100010100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10100010101000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10100010101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10100010101010) && ({row_reg, col_reg}<14'b10100010101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100010101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10100010101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10100010101110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10100010101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10100010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10100010110001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10100010110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10100010110011) && ({row_reg, col_reg}<14'b10100010110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10100010110111) && ({row_reg, col_reg}<14'b10100010111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10100010111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10100010111100) && ({row_reg, col_reg}<14'b10100011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10100011000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=14'b10100011000010) && ({row_reg, col_reg}<14'b10100011000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10100011000110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=14'b10100011000111) && ({row_reg, col_reg}<14'b10100011001010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=14'b10100011001010) && ({row_reg, col_reg}<14'b10100011001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10100011001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10100011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10100011001111)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b10100011010000) && ({row_reg, col_reg}<14'b10100100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100100011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10100100011001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==14'b10100100011010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10100100011011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b10100100011100)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}>=14'b10100100011101) && ({row_reg, col_reg}<14'b10100100100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10100100100001) && ({row_reg, col_reg}<14'b10100100100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10100100100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10100100100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10100100100101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10100100100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b10100100100111) && ({row_reg, col_reg}<14'b10100100101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10100100101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b10100100101011) && ({row_reg, col_reg}<14'b10100100101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10100100101101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10100100101110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10100100101111) && ({row_reg, col_reg}<14'b10100100110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10100100110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10100100110010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10100100110011) && ({row_reg, col_reg}<14'b10100100110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10100100110111) && ({row_reg, col_reg}<14'b10100100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10100100111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10100100111100) && ({row_reg, col_reg}<14'b10100101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10100101000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==14'b10100101000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=14'b10100101000011) && ({row_reg, col_reg}<14'b10100101000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b10100101000101) && ({row_reg, col_reg}<14'b10100101000111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=14'b10100101000111) && ({row_reg, col_reg}<14'b10100101001001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10100101001001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=14'b10100101001010) && ({row_reg, col_reg}<14'b10100101001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b10100101001100) && ({row_reg, col_reg}<14'b10100101001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10100101001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10100101001111)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b10100101010000) && ({row_reg, col_reg}<14'b10100110010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100110010111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b10100110011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b10100110011001) && ({row_reg, col_reg}<14'b10100110011011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b10100110011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b10100110011100) && ({row_reg, col_reg}<14'b10100110100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10100110100000) && ({row_reg, col_reg}<14'b10100110100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10100110100010) && ({row_reg, col_reg}<14'b10100110100100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10100110100100) && ({row_reg, col_reg}<14'b10100110100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10100110100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10100110100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b10100110101000) && ({row_reg, col_reg}<14'b10100110101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10100110101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10100110101011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10100110101100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10100110101101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10100110101110) && ({row_reg, col_reg}<14'b10100110110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10100110110000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10100110110001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10100110110010) && ({row_reg, col_reg}<14'b10100110110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10100110110111) && ({row_reg, col_reg}<14'b10100110111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10100110111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10100110111100) && ({row_reg, col_reg}<14'b10100111000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10100111000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==14'b10100111000010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=14'b10100111000011) && ({row_reg, col_reg}<14'b10100111001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b10100111001010) && ({row_reg, col_reg}<14'b10100111001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=14'b10100111001100) && ({row_reg, col_reg}<14'b10100111001111)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=14'b10100111001111) && ({row_reg, col_reg}<14'b10101000010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101000010111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b10101000011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b10101000011001) && ({row_reg, col_reg}<14'b10101000011100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=14'b10101000011100) && ({row_reg, col_reg}<14'b10101000100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10101000100000) && ({row_reg, col_reg}<14'b10101000100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10101000100010) && ({row_reg, col_reg}<14'b10101000100100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10101000100100) && ({row_reg, col_reg}<14'b10101000100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10101000100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10101000100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b10101000101000) && ({row_reg, col_reg}<14'b10101000101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10101000101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10101000101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b10101000101100) && ({row_reg, col_reg}<14'b10101000101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10101000101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10101000110000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10101000110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10101000110010) && ({row_reg, col_reg}<14'b10101000110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10101000110110) && ({row_reg, col_reg}<14'b10101000111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10101000111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10101000111100) && ({row_reg, col_reg}<14'b10101001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10101001000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=14'b10101001000010) && ({row_reg, col_reg}<14'b10101001001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10101001001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=14'b10101001001011) && ({row_reg, col_reg}<14'b10101001001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10101001001110)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b10101001001111) && ({row_reg, col_reg}<14'b10101010010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10101010010110) && ({row_reg, col_reg}<14'b10101010011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10101010011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10101010011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10101010011010) && ({row_reg, col_reg}<14'b10101010100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10101010100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10101010100001) && ({row_reg, col_reg}<14'b10101010100100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10101010100100) && ({row_reg, col_reg}<14'b10101010100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10101010100110) && ({row_reg, col_reg}<14'b10101010101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10101010101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10101010101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10101010101011) && ({row_reg, col_reg}<14'b10101010101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10101010101101) && ({row_reg, col_reg}<14'b10101010101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10101010101111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10101010110000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10101010110001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10101010110010) && ({row_reg, col_reg}<14'b10101010110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10101010110110) && ({row_reg, col_reg}<14'b10101010111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10101010111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10101010111011) && ({row_reg, col_reg}<14'b10101011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10101011000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==14'b10101011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b10101011000010) && ({row_reg, col_reg}<14'b10101011000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b10101011000110) && ({row_reg, col_reg}<14'b10101011001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=14'b10101011001000) && ({row_reg, col_reg}<14'b10101011001010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b10101011001010) && ({row_reg, col_reg}<14'b10101011001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b10101011001100) && ({row_reg, col_reg}<14'b10101011001111)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b10101011001111) && ({row_reg, col_reg}<14'b10101100010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10101100010110) && ({row_reg, col_reg}<14'b10101100011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10101100011001) && ({row_reg, col_reg}<14'b10101100100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10101100100000) && ({row_reg, col_reg}<14'b10101100100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10101100100111) && ({row_reg, col_reg}<14'b10101100101001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10101100101001) && ({row_reg, col_reg}<14'b10101100101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10101100101011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10101100101100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b10101100101101) && ({row_reg, col_reg}<14'b10101100110000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10101100110000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10101100110001) && ({row_reg, col_reg}<14'b10101100110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10101100110110) && ({row_reg, col_reg}<14'b10101100111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10101100111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10101100111011) && ({row_reg, col_reg}<14'b10101101000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10101101000000) && ({row_reg, col_reg}<14'b10101101000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b10101101000111) && ({row_reg, col_reg}<14'b10101101001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=14'b10101101001010) && ({row_reg, col_reg}<14'b10101101001100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b10101101001100) && ({row_reg, col_reg}<14'b10101101001111)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b10101101001111) && ({row_reg, col_reg}<14'b10101110010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101110010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10101110010110) && ({row_reg, col_reg}<14'b10101110011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10101110011111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10101110100000) && ({row_reg, col_reg}<14'b10101110100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10101110100011) && ({row_reg, col_reg}<14'b10101110100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10101110100110) && ({row_reg, col_reg}<14'b10101110101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10101110101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b10101110101011) && ({row_reg, col_reg}<14'b10101110101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10101110101110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10101110101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10101110110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10101110110001) && ({row_reg, col_reg}<14'b10101110110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10101110110110) && ({row_reg, col_reg}<14'b10101110111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10101110111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10101110111011) && ({row_reg, col_reg}<14'b10101110111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10101110111111) && ({row_reg, col_reg}<14'b10101111000010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b10101111000010) && ({row_reg, col_reg}<14'b10101111000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10101111000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10101111000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b10101111000111) && ({row_reg, col_reg}<14'b10101111001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10101111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10101111001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=14'b10101111001011) && ({row_reg, col_reg}<14'b10101111001101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10101111001101)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b10101111001110) && ({row_reg, col_reg}<14'b10110000010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10110000010101) && ({row_reg, col_reg}<14'b10110000011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10110000011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110000011001) && ({row_reg, col_reg}<14'b10110000011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10110000011110) && ({row_reg, col_reg}<14'b10110000100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10110000100000) && ({row_reg, col_reg}<14'b10110000100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10110000100101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10110000100110) && ({row_reg, col_reg}<14'b10110000101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10110000101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b10110000101011) && ({row_reg, col_reg}<14'b10110000101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10110000101101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10110000101110) && ({row_reg, col_reg}<14'b10110000110000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10110000110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10110000110001) && ({row_reg, col_reg}<14'b10110000110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10110000110101) && ({row_reg, col_reg}<14'b10110000111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10110000111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10110000111010) && ({row_reg, col_reg}<14'b10110000111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10110000111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10110001000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10110001000001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=14'b10110001000010) && ({row_reg, col_reg}<14'b10110001000100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10110001000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b10110001000101) && ({row_reg, col_reg}<14'b10110001000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10110001000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10110001001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=14'b10110001001001) && ({row_reg, col_reg}<14'b10110001001011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10110001001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==14'b10110001001100)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=14'b10110001001101) && ({row_reg, col_reg}<14'b10110010010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10110010010101) && ({row_reg, col_reg}<14'b10110010011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10110010011000) && ({row_reg, col_reg}<14'b10110010011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110010011010) && ({row_reg, col_reg}<14'b10110010011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10110010011110) && ({row_reg, col_reg}<14'b10110010100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10110010100000) && ({row_reg, col_reg}<14'b10110010100100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10110010100100) && ({row_reg, col_reg}<14'b10110010100111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10110010100111) && ({row_reg, col_reg}<14'b10110010101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10110010101101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10110010101110) && ({row_reg, col_reg}<14'b10110010110000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10110010110000) && ({row_reg, col_reg}<14'b10110010110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10110010110101) && ({row_reg, col_reg}<14'b10110010111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10110010111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10110010111010) && ({row_reg, col_reg}<14'b10110010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10110010111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10110011000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10110011000001)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==14'b10110011000010)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==14'b10110011000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10110011000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10110011000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b10110011000110) && ({row_reg, col_reg}<14'b10110011001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10110011001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b10110011001010) && ({row_reg, col_reg}<14'b10110011001101)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b10110011001101) && ({row_reg, col_reg}<14'b10110100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10110100010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110100010101) && ({row_reg, col_reg}<14'b10110100011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10110100011000) && ({row_reg, col_reg}<14'b10110100011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110100011011) && ({row_reg, col_reg}<14'b10110100011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10110100011110) && ({row_reg, col_reg}<14'b10110100100001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10110100100001) && ({row_reg, col_reg}<14'b10110100100100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10110100100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10110100100101) && ({row_reg, col_reg}<14'b10110100101100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b10110100101100) && ({row_reg, col_reg}<14'b10110100101110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10110100101110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10110100101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10110100110000) && ({row_reg, col_reg}<14'b10110100110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10110100110101) && ({row_reg, col_reg}<14'b10110100111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10110100111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10110100111010) && ({row_reg, col_reg}<14'b10110100111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10110100111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10110101000000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=14'b10110101000001) && ({row_reg, col_reg}<14'b10110101000011)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==14'b10110101000011)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==14'b10110101000100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b10110101000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10110101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b10110101000111) && ({row_reg, col_reg}<14'b10110101001010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=14'b10110101001010) && ({row_reg, col_reg}<14'b10110101001100)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b10110101001100) && ({row_reg, col_reg}<14'b10110110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10110110010100) && ({row_reg, col_reg}<14'b10110110010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10110110010111) && ({row_reg, col_reg}<14'b10110110011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110110011011) && ({row_reg, col_reg}<14'b10110110011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10110110011110) && ({row_reg, col_reg}<14'b10110110100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10110110100000) && ({row_reg, col_reg}<14'b10110110100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10110110100011) && ({row_reg, col_reg}<14'b10110110100101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10110110100101) && ({row_reg, col_reg}<14'b10110110101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10110110101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b10110110101001) && ({row_reg, col_reg}<14'b10110110101100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10110110101100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10110110101101) && ({row_reg, col_reg}<14'b10110110101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10110110101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10110110110000) && ({row_reg, col_reg}<14'b10110110110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10110110110101) && ({row_reg, col_reg}<14'b10110110111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10110110111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10110110111010) && ({row_reg, col_reg}<14'b10110110111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10110110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10110110111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10110111000000)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}>=14'b10110111000001) && ({row_reg, col_reg}<14'b10110111000011)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==14'b10110111000011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b10110111000100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=14'b10110111000101) && ({row_reg, col_reg}<14'b10110111001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10110111001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10110111001010)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b10110111001011) && ({row_reg, col_reg}<14'b10111000010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111000010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10111000010100) && ({row_reg, col_reg}<14'b10111000010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10111000010111) && ({row_reg, col_reg}<14'b10111000011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10111000011011) && ({row_reg, col_reg}<14'b10111000011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10111000011110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10111000011111) && ({row_reg, col_reg}<14'b10111000100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10111000100011) && ({row_reg, col_reg}<14'b10111000100101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10111000100101) && ({row_reg, col_reg}<14'b10111000100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b10111000100111) && ({row_reg, col_reg}<14'b10111000101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b10111000101010) && ({row_reg, col_reg}<14'b10111000101100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10111000101100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10111000101101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10111000101110) && ({row_reg, col_reg}<14'b10111000110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10111000110000) && ({row_reg, col_reg}<14'b10111000110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10111000110100) && ({row_reg, col_reg}<14'b10111000111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10111000111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10111000111111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10111001000000)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==14'b10111001000001)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==14'b10111001000010)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==14'b10111001000011)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==14'b10111001000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b10111001000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10111001000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10111001000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10111001001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10111001001001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10111001001010)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b10111001001011) && ({row_reg, col_reg}<14'b10111010010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10111010010011) && ({row_reg, col_reg}<14'b10111010010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10111010010111) && ({row_reg, col_reg}<14'b10111010011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10111010011011) && ({row_reg, col_reg}<14'b10111010011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10111010011110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10111010011111) && ({row_reg, col_reg}<14'b10111010100010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10111010100010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10111010100011) && ({row_reg, col_reg}<14'b10111010100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b10111010100110) && ({row_reg, col_reg}<14'b10111010101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10111010101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b10111010101011) && ({row_reg, col_reg}<14'b10111010101101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10111010101101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10111010101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10111010101111) && ({row_reg, col_reg}<14'b10111010110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10111010110100) && ({row_reg, col_reg}<14'b10111010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10111010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10111010111001) && ({row_reg, col_reg}<14'b10111010111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10111010111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10111010111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10111011000000)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}>=14'b10111011000001) && ({row_reg, col_reg}<14'b10111011000011)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==14'b10111011000011)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==14'b10111011000100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b10111011000101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=14'b10111011000110) && ({row_reg, col_reg}<14'b10111011001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10111011001001)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=14'b10111011001010) && ({row_reg, col_reg}<14'b10111100010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10111100010011) && ({row_reg, col_reg}<14'b10111100010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10111100010110) && ({row_reg, col_reg}<14'b10111100011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10111100011010) && ({row_reg, col_reg}<14'b10111100011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10111100011101) && ({row_reg, col_reg}<14'b10111100011111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10111100011111) && ({row_reg, col_reg}<14'b10111100100010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10111100100010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10111100100011) && ({row_reg, col_reg}<14'b10111100100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b10111100100110) && ({row_reg, col_reg}<14'b10111100101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10111100101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10111100101011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10111100101100) && ({row_reg, col_reg}<14'b10111100101110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10111100101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10111100101111) && ({row_reg, col_reg}<14'b10111100110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10111100110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10111100110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10111100110110) && ({row_reg, col_reg}<14'b10111100111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10111100111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10111100111001) && ({row_reg, col_reg}<14'b10111100111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10111100111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10111100111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=14'b10111101000000) && ({row_reg, col_reg}<14'b10111101000010)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}>=14'b10111101000010) && ({row_reg, col_reg}<14'b10111101000100)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==14'b10111101000100)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==14'b10111101000101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b10111101000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b10111101000111) && ({row_reg, col_reg}<14'b10111101001010)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=14'b10111101001010) && ({row_reg, col_reg}<14'b10111110010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10111110010010) && ({row_reg, col_reg}<14'b10111110010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10111110010110) && ({row_reg, col_reg}<14'b10111110011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10111110011001) && ({row_reg, col_reg}<14'b10111110011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10111110011110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10111110011111) && ({row_reg, col_reg}<14'b10111110100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10111110100001) && ({row_reg, col_reg}<14'b10111110100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10111110100011) && ({row_reg, col_reg}<14'b10111110100101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b10111110100101) && ({row_reg, col_reg}<14'b10111110100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10111110100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b10111110101000) && ({row_reg, col_reg}<14'b10111110101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10111110101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10111110101011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10111110101100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10111110101101) && ({row_reg, col_reg}<14'b10111110101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10111110101111) && ({row_reg, col_reg}<14'b10111110110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10111110110100) && ({row_reg, col_reg}<14'b10111110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10111110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10111110111001) && ({row_reg, col_reg}<14'b10111110111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10111110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10111110111111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b10111111000000)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}>=14'b10111111000001) && ({row_reg, col_reg}<14'b10111111000011)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==14'b10111111000011)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b10111111000100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b10111111000101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b10111111000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10111111000111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b10111111001000)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b10111111001001) && ({row_reg, col_reg}<14'b11000000010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b11000000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11000000010010) && ({row_reg, col_reg}<14'b11000000010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b11000000010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11000000010110) && ({row_reg, col_reg}<14'b11000000011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b11000000011110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11000000011111) && ({row_reg, col_reg}<14'b11000000100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11000000100001) && ({row_reg, col_reg}<14'b11000000100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b11000000100011) && ({row_reg, col_reg}<14'b11000000100101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b11000000100101) && ({row_reg, col_reg}<14'b11000000100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b11000000100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b11000000101000) && ({row_reg, col_reg}<14'b11000000101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b11000000101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b11000000101011) && ({row_reg, col_reg}<14'b11000000101101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11000000101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11000000101110) && ({row_reg, col_reg}<14'b11000000110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11000000110100) && ({row_reg, col_reg}<14'b11000000111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11000000111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11000000111001) && ({row_reg, col_reg}<14'b11000000111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11000000111101) && ({row_reg, col_reg}<14'b11000000111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b11000000111111) && ({row_reg, col_reg}<14'b11000001000010)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==14'b11000001000010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b11000001000011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b11000001000100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b11000001000101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b11000001000110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11000001000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b11000001001000)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b11000001001001) && ({row_reg, col_reg}<14'b11000010010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b11000010010000) && ({row_reg, col_reg}<14'b11000010010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11000010010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11000010010100) && ({row_reg, col_reg}<14'b11000010011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11000010011010) && ({row_reg, col_reg}<14'b11000010100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11000010100000) && ({row_reg, col_reg}<14'b11000010100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11000010100011) && ({row_reg, col_reg}<14'b11000010100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11000010100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11000010100111) && ({row_reg, col_reg}<14'b11000010101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11000010101010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b11000010101011) && ({row_reg, col_reg}<14'b11000010101101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11000010101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11000010101110) && ({row_reg, col_reg}<14'b11000010110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b11000010110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11000010110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b11000010110101) && ({row_reg, col_reg}<14'b11000010110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11000010110111) && ({row_reg, col_reg}<14'b11000010111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11000010111001) && ({row_reg, col_reg}<14'b11000010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11000010111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b11000010111110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=14'b11000010111111) && ({row_reg, col_reg}<14'b11000011000001)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==14'b11000011000001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b11000011000010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b11000011000011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b11000011000100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=14'b11000011000101) && ({row_reg, col_reg}<14'b11000011000111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11000011000111)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}>=14'b11000011001000) && ({row_reg, col_reg}<14'b11000100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b11000100001110) && ({row_reg, col_reg}<14'b11000100010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11000100010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b11000100010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11000100010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11000100010110) && ({row_reg, col_reg}<14'b11000100011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11000100011000) && ({row_reg, col_reg}<14'b11000100011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11000100011111) && ({row_reg, col_reg}<14'b11000100100101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11000100100101) && ({row_reg, col_reg}<14'b11000100101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11000100101010) && ({row_reg, col_reg}<14'b11000100101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b11000100101101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11000100101110) && ({row_reg, col_reg}<14'b11000100110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b11000100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11000100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b11000100110101) && ({row_reg, col_reg}<14'b11000100110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11000100110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11000100111000) && ({row_reg, col_reg}<14'b11000100111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11000100111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b11000100111110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11000100111111)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}>=14'b11000101000000) && ({row_reg, col_reg}<14'b11000101000010)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b11000101000010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b11000101000011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=14'b11000101000100) && ({row_reg, col_reg}<14'b11000101000110)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}>=14'b11000101000110) && ({row_reg, col_reg}<14'b11000110001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b11000110001101) && ({row_reg, col_reg}<14'b11000110001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11000110001111) && ({row_reg, col_reg}<14'b11000110011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11000110011101) && ({row_reg, col_reg}<14'b11000110100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11000110100100) && ({row_reg, col_reg}<14'b11000110101101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11000110101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11000110101110) && ({row_reg, col_reg}<14'b11000110110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11000110110011) && ({row_reg, col_reg}<14'b11000110110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11000110110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11000110111000) && ({row_reg, col_reg}<14'b11000110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11000110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b11000110111110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b11000110111111) && ({row_reg, col_reg}<14'b11000111000001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==14'b11000111000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b11000111000010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b11000111000011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b11000111000100)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}>=14'b11000111000101) && ({row_reg, col_reg}<14'b11001000001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b11001000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11001000001101) && ({row_reg, col_reg}<14'b11001000011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11001000011011) && ({row_reg, col_reg}<14'b11001000100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11001000100100) && ({row_reg, col_reg}<14'b11001000101110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11001000101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11001000101111) && ({row_reg, col_reg}<14'b11001000110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11001000110011) && ({row_reg, col_reg}<14'b11001000110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11001000110110) && ({row_reg, col_reg}<14'b11001000111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11001000111000) && ({row_reg, col_reg}<14'b11001000111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11001000111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b11001000111110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b11001000111111) && ({row_reg, col_reg}<14'b11001001000001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b11001001000001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b11001001000010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=14'b11001001000011) && ({row_reg, col_reg}<14'b11001001000101)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}>=14'b11001001000101) && ({row_reg, col_reg}<14'b11001010001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b11001010001011) && ({row_reg, col_reg}<14'b11001010001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11001010001101) && ({row_reg, col_reg}<14'b11001010011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11001010011100) && ({row_reg, col_reg}<14'b11001010100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11001010100100) && ({row_reg, col_reg}<14'b11001010101110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11001010101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11001010101111) && ({row_reg, col_reg}<14'b11001010110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11001010110001) && ({row_reg, col_reg}<14'b11001010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11001010110110) && ({row_reg, col_reg}<14'b11001010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11001010111000) && ({row_reg, col_reg}<14'b11001010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11001010111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==14'b11001010111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b11001010111110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b11001010111111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b11001011000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b11001011000001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=14'b11001011000010) && ({row_reg, col_reg}<14'b11001011000101)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}>=14'b11001011000101) && ({row_reg, col_reg}<14'b11001100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b11001100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11001100001100) && ({row_reg, col_reg}<14'b11001100011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11001100011011) && ({row_reg, col_reg}<14'b11001100100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11001100100100) && ({row_reg, col_reg}<14'b11001100101110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11001100101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11001100101111) && ({row_reg, col_reg}<14'b11001100110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11001100110001) && ({row_reg, col_reg}<14'b11001100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11001100110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11001100110111) && ({row_reg, col_reg}<14'b11001100111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11001100111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b11001100111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=14'b11001100111110) && ({row_reg, col_reg}<14'b11001101000001)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=14'b11001101000001) && ({row_reg, col_reg}<14'b11001101000100)) color_data = 12'b001100100001;

		if(({row_reg, col_reg}>=14'b11001101000100) && ({row_reg, col_reg}<14'b11001110001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b11001110001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11001110001011) && ({row_reg, col_reg}<14'b11001110011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11001110011010) && ({row_reg, col_reg}<14'b11001110100001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b11001110100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11001110100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11001110100011) && ({row_reg, col_reg}<14'b11001110100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11001110100101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b11001110100110) && ({row_reg, col_reg}<14'b11001110101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11001110101011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11001110101100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11001110101101) && ({row_reg, col_reg}<14'b11001110101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11001110101111) && ({row_reg, col_reg}<14'b11001110110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11001110110010) && ({row_reg, col_reg}<14'b11001110110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11001110110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11001110110111) && ({row_reg, col_reg}<14'b11001110111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11001110111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b11001110111101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b11001110111110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=14'b11001110111111) && ({row_reg, col_reg}<14'b11001111000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11001111000011)) color_data = 12'b001000100000;

		if(({row_reg, col_reg}>=14'b11001111000100) && ({row_reg, col_reg}<14'b11010000001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b11010000001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11010000001011) && ({row_reg, col_reg}<14'b11010000011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11010000011001) && ({row_reg, col_reg}<14'b11010000100001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11010000100001) && ({row_reg, col_reg}<14'b11010000100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11010000100110) && ({row_reg, col_reg}<14'b11010000101001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b11010000101001) && ({row_reg, col_reg}<14'b11010000101101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11010000101101) && ({row_reg, col_reg}<14'b11010000101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11010000101111) && ({row_reg, col_reg}<14'b11010000110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11010000110011) && ({row_reg, col_reg}<14'b11010000111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11010000111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b11010000111101) && ({row_reg, col_reg}<14'b11010001000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11010001000011)) color_data = 12'b001000100000;

		if(({row_reg, col_reg}>=14'b11010001000100) && ({row_reg, col_reg}<14'b11010010001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b11010010001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11010010001010) && ({row_reg, col_reg}<14'b11010010011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11010010011001) && ({row_reg, col_reg}<14'b11010010100001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11010010100001) && ({row_reg, col_reg}<14'b11010010100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11010010100110) && ({row_reg, col_reg}<14'b11010010101100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11010010101100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11010010101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11010010101110) && ({row_reg, col_reg}<14'b11010010110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11010010110011) && ({row_reg, col_reg}<14'b11010010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11010010111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b11010010111101) && ({row_reg, col_reg}<14'b11010011000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11010011000010)) color_data = 12'b001000100000;

		if(({row_reg, col_reg}>=14'b11010011000011) && ({row_reg, col_reg}<14'b11010100001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b11010100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11010100001010) && ({row_reg, col_reg}<14'b11010100011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11010100011000) && ({row_reg, col_reg}<14'b11010100100001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11010100100001) && ({row_reg, col_reg}<14'b11010100100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11010100100110) && ({row_reg, col_reg}<14'b11010100101011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b11010100101011) && ({row_reg, col_reg}<14'b11010100101101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11010100101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11010100101110) && ({row_reg, col_reg}<14'b11010100110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11010100110100) && ({row_reg, col_reg}<14'b11010100111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11010100111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b11010100111101) && ({row_reg, col_reg}<14'b11010101000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11010101000010)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}>=14'b11010101000011) && ({row_reg, col_reg}<14'b11010110001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b11010110001001) && ({row_reg, col_reg}<14'b11010110011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11010110011000) && ({row_reg, col_reg}<14'b11010110100001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11010110100001) && ({row_reg, col_reg}<14'b11010110101000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11010110101000) && ({row_reg, col_reg}<14'b11010110101011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b11010110101011) && ({row_reg, col_reg}<14'b11010110101101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11010110101101) && ({row_reg, col_reg}<14'b11010110110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11010110110101) && ({row_reg, col_reg}<14'b11010110111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11010110111011) && ({row_reg, col_reg}<14'b11010110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b11010110111101) && ({row_reg, col_reg}<14'b11010111000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11010111000001)) color_data = 12'b001000100000;

		if(({row_reg, col_reg}>=14'b11010111000010) && ({row_reg, col_reg}<14'b11011000001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b11011000001000) && ({row_reg, col_reg}<14'b11011000010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11011000010111) && ({row_reg, col_reg}<14'b11011000100001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11011000100001) && ({row_reg, col_reg}<14'b11011000100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11011000100011) && ({row_reg, col_reg}<14'b11011000100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11011000100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11011000100111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b11011000101000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11011000101001) && ({row_reg, col_reg}<14'b11011000101011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11011000101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11011000101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11011000101101) && ({row_reg, col_reg}<14'b11011000110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11011000110101) && ({row_reg, col_reg}<14'b11011000111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11011000111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b11011000111011) && ({row_reg, col_reg}<14'b11011000111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b11011000111101) && ({row_reg, col_reg}<14'b11011001000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b11011001000000) && ({row_reg, col_reg}<14'b11011001000010)) color_data = 12'b001000100000;

		if(({row_reg, col_reg}>=14'b11011001000010) && ({row_reg, col_reg}<14'b11011010001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b11011010001000) && ({row_reg, col_reg}<14'b11011010010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11011010010101) && ({row_reg, col_reg}<14'b11011010011001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b11011010011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11011010011010) && ({row_reg, col_reg}<14'b11011010100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11011010100000) && ({row_reg, col_reg}<14'b11011010100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11011010100011) && ({row_reg, col_reg}<14'b11011010100111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11011010100111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11011010101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b11011010101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11011010101010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11011010101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11011010101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11011010101101) && ({row_reg, col_reg}<14'b11011010110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11011010110110) && ({row_reg, col_reg}<14'b11011010111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11011010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b11011010111011) && ({row_reg, col_reg}<14'b11011010111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b11011010111101) && ({row_reg, col_reg}<14'b11011011000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11011011000000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b11011011000001)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}>=14'b11011011000010) && ({row_reg, col_reg}<14'b11011100001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b11011100001000) && ({row_reg, col_reg}<14'b11011100010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11011100010100) && ({row_reg, col_reg}<14'b11011100100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11011100100000) && ({row_reg, col_reg}<14'b11011100100010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11011100100010) && ({row_reg, col_reg}<14'b11011100101000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b11011100101000) && ({row_reg, col_reg}<14'b11011100101100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11011100101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11011100101101) && ({row_reg, col_reg}<14'b11011100110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11011100110111) && ({row_reg, col_reg}<14'b11011100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11011100111011) && ({row_reg, col_reg}<14'b11011100111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=14'b11011100111101) && ({row_reg, col_reg}<14'b11011101000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11011101000000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b11011101000001)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}>=14'b11011101000010) && ({row_reg, col_reg}<14'b11011110000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b11011110000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11011110001000) && ({row_reg, col_reg}<14'b11011110010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11011110010101) && ({row_reg, col_reg}<14'b11011110011111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11011110011111) && ({row_reg, col_reg}<14'b11011110100010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11011110100010) && ({row_reg, col_reg}<14'b11011110101001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b11011110101001) && ({row_reg, col_reg}<14'b11011110101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11011110101011) && ({row_reg, col_reg}<14'b11011110101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11011110101101) && ({row_reg, col_reg}<14'b11011110110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11011110110111) && ({row_reg, col_reg}<14'b11011110111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11011110111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b11011110111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=14'b11011110111101) && ({row_reg, col_reg}<14'b11011110111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b11011110111111) && ({row_reg, col_reg}<14'b11011111000001)) color_data = 12'b001000100000;

		if(({row_reg, col_reg}>=14'b11011111000001) && ({row_reg, col_reg}<14'b11100000000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b11100000000111) && ({row_reg, col_reg}<14'b11100000010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b11100000010100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11100000010101) && ({row_reg, col_reg}<14'b11100000010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11100000010111) && ({row_reg, col_reg}<14'b11100000011111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11100000011111) && ({row_reg, col_reg}<14'b11100000100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11100000100001) && ({row_reg, col_reg}<14'b11100000101010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b11100000101010) && ({row_reg, col_reg}<14'b11100000101100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11100000101100) && ({row_reg, col_reg}<14'b11100000111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11100000111000) && ({row_reg, col_reg}<14'b11100000111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11100000111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b11100000111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=14'b11100000111101) && ({row_reg, col_reg}<14'b11100000111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11100000111111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b11100001000000)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}>=14'b11100001000001) && ({row_reg, col_reg}<14'b11100010000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b11100010000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11100010000111) && ({row_reg, col_reg}<14'b11100010010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11100010010110) && ({row_reg, col_reg}<14'b11100010011111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11100010011111) && ({row_reg, col_reg}<14'b11100010100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11100010100001) && ({row_reg, col_reg}<14'b11100010101010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11100010101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11100010101011) && ({row_reg, col_reg}<14'b11100010101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11100010101101) && ({row_reg, col_reg}<14'b11100010101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b11100010101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11100010110000) && ({row_reg, col_reg}<14'b11100010110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b11100010110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11100010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11100010111001) && ({row_reg, col_reg}<14'b11100010111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11100010111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==14'b11100010111100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=14'b11100010111101) && ({row_reg, col_reg}<14'b11100010111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11100010111111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b11100011000000)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}>=14'b11100011000001) && ({row_reg, col_reg}<14'b11100100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b11100100000110) && ({row_reg, col_reg}<14'b11100100010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11100100010110) && ({row_reg, col_reg}<14'b11100100011101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11100100011101) && ({row_reg, col_reg}<14'b11100100100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11100100100001) && ({row_reg, col_reg}<14'b11100100101001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11100100101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b11100100101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11100100101011) && ({row_reg, col_reg}<14'b11100100111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11100100111000) && ({row_reg, col_reg}<14'b11100100111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11100100111100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b11100100111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11100100111110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b11100100111111)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}>=14'b11100101000000) && ({row_reg, col_reg}<14'b11100110000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b11100110000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11100110000110) && ({row_reg, col_reg}<14'b11100110010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11100110010111) && ({row_reg, col_reg}<14'b11100110011101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11100110011101) && ({row_reg, col_reg}<14'b11100110100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11100110100001) && ({row_reg, col_reg}<14'b11100110101001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11100110101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b11100110101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11100110101011) && ({row_reg, col_reg}<14'b11100110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11100110111000) && ({row_reg, col_reg}<14'b11100110111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11100110111100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b11100110111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11100110111110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b11100110111111)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=14'b11100111000000) && ({row_reg, col_reg}<14'b11101000000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b11101000000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11101000000110) && ({row_reg, col_reg}<14'b11101000010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11101000010111) && ({row_reg, col_reg}<14'b11101000011100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11101000011100) && ({row_reg, col_reg}<14'b11101000100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11101000100000) && ({row_reg, col_reg}<14'b11101000101001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11101000101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b11101000101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11101000101011) && ({row_reg, col_reg}<14'b11101000111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11101000111000) && ({row_reg, col_reg}<14'b11101000111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11101000111100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b11101000111101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11101000111110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b11101000111111)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=14'b11101001000000) && ({row_reg, col_reg}<14'b11101010000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b11101010000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11101010000110) && ({row_reg, col_reg}<14'b11101010010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11101010010110) && ({row_reg, col_reg}<14'b11101010011010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11101010011010) && ({row_reg, col_reg}<14'b11101010100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11101010100001) && ({row_reg, col_reg}<14'b11101010101000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11101010101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b11101010101001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11101010101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b11101010101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b11101010101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11101010101101) && ({row_reg, col_reg}<14'b11101010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11101010111000) && ({row_reg, col_reg}<14'b11101010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11101010111100) && ({row_reg, col_reg}<14'b11101010111110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b11101010111110)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}>=14'b11101010111111) && ({row_reg, col_reg}<14'b11101100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b11101100000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11101100000101) && ({row_reg, col_reg}<14'b11101100010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11101100010110) && ({row_reg, col_reg}<14'b11101100011001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11101100011001) && ({row_reg, col_reg}<14'b11101100100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11101100100000) && ({row_reg, col_reg}<14'b11101100101000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11101100101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b11101100101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11101100101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b11101100101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b11101100101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11101100101101) && ({row_reg, col_reg}<14'b11101100111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11101100111000) && ({row_reg, col_reg}<14'b11101100111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11101100111100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11101100111101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b11101100111110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=14'b11101100111111) && ({row_reg, col_reg}<14'b11101110000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b11101110000011) && ({row_reg, col_reg}<14'b11101110000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11101110000101) && ({row_reg, col_reg}<14'b11101110010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11101110010110) && ({row_reg, col_reg}<14'b11101110011001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11101110011001) && ({row_reg, col_reg}<14'b11101110011111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11101110011111) && ({row_reg, col_reg}<14'b11101110101000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11101110101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b11101110101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11101110101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11101110101011) && ({row_reg, col_reg}<14'b11101110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11101110111000) && ({row_reg, col_reg}<14'b11101110111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11101110111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==14'b11101110111100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11101110111101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b11101110111110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=14'b11101110111111) && ({row_reg, col_reg}<14'b11110000000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b11110000000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11110000000100) && ({row_reg, col_reg}<14'b11110000010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11110000010101) && ({row_reg, col_reg}<14'b11110000011001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11110000011001) && ({row_reg, col_reg}<14'b11110000100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11110000100000) && ({row_reg, col_reg}<14'b11110000101000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11110000101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b11110000101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11110000101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b11110000101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11110000101100) && ({row_reg, col_reg}<14'b11110000101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11110000101110) && ({row_reg, col_reg}<14'b11110000111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11110000111000) && ({row_reg, col_reg}<14'b11110000111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11110000111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b11110000111100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==14'b11110000111101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b11110000111110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=14'b11110000111111) && ({row_reg, col_reg}<14'b11110010000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b11110010000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11110010000100) && ({row_reg, col_reg}<14'b11110010010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11110010010110) && ({row_reg, col_reg}<14'b11110010011001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11110010011001) && ({row_reg, col_reg}<14'b11110010011111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11110010011111) && ({row_reg, col_reg}<14'b11110010101001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b11110010101001) && ({row_reg, col_reg}<14'b11110010101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b11110010101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b11110010101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11110010101110) && ({row_reg, col_reg}<14'b11110010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11110010111000) && ({row_reg, col_reg}<14'b11110010111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11110010111011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b11110010111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b11110010111101)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=14'b11110010111110) && ({row_reg, col_reg}<14'b11110100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b11110100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11110100000011) && ({row_reg, col_reg}<14'b11110100010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11110100010101) && ({row_reg, col_reg}<14'b11110100011001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11110100011001) && ({row_reg, col_reg}<14'b11110100011110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11110100011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11110100011111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b11110100100000) && ({row_reg, col_reg}<14'b11110100101000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11110100101000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11110100101001) && ({row_reg, col_reg}<14'b11110100101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b11110100101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b11110100101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11110100110000) && ({row_reg, col_reg}<14'b11110100111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11110100111000) && ({row_reg, col_reg}<14'b11110100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11110100111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==14'b11110100111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b11110100111101)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}>=14'b11110100111110) && ({row_reg, col_reg}<14'b11110110000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b11110110000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11110110000011) && ({row_reg, col_reg}<14'b11110110010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11110110010101) && ({row_reg, col_reg}<14'b11110110011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11110110011000) && ({row_reg, col_reg}<14'b11110110011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11110110011101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b11110110011110) && ({row_reg, col_reg}<14'b11110110100000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b11110110100000) && ({row_reg, col_reg}<14'b11110110100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b11110110100110) && ({row_reg, col_reg}<14'b11110110101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b11110110101000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11110110101001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b11110110101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11110110101011) && ({row_reg, col_reg}<14'b11110110101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b11110110101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b11110110101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11110110110000) && ({row_reg, col_reg}<14'b11110110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11110110111000) && ({row_reg, col_reg}<14'b11110110111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11110110111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==14'b11110110111100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b11110110111101)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b11110110111110) && ({row_reg, col_reg}<14'b11111000000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b11111000000001) && ({row_reg, col_reg}<14'b11111000000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11111000000011) && ({row_reg, col_reg}<14'b11111000010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11111000010011) && ({row_reg, col_reg}<14'b11111000011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11111000011000) && ({row_reg, col_reg}<14'b11111000011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11111000011101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11111000011110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b11111000011111) && ({row_reg, col_reg}<14'b11111000100001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11111000100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b11111000100010) && ({row_reg, col_reg}<14'b11111000100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b11111000100100) && ({row_reg, col_reg}<14'b11111000100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b11111000100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11111000100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b11111000101000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11111000101001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11111000101010) && ({row_reg, col_reg}<14'b11111000101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b11111000101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11111000101101) && ({row_reg, col_reg}<14'b11111000111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11111000111000) && ({row_reg, col_reg}<14'b11111000111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b11111000111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b11111000111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==14'b11111000111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==14'b11111000111101)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b11111000111110) && ({row_reg, col_reg}<14'b11111010000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b11111010000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11111010000010) && ({row_reg, col_reg}<14'b11111010010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11111010010011) && ({row_reg, col_reg}<14'b11111010011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11111010011000) && ({row_reg, col_reg}<14'b11111010011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11111010011101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11111010011110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b11111010011111) && ({row_reg, col_reg}<14'b11111010100111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11111010100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b11111010101000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11111010101001) && ({row_reg, col_reg}<14'b11111010101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11111010101101) && ({row_reg, col_reg}<14'b11111010101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b11111010101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11111010110000) && ({row_reg, col_reg}<14'b11111010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11111010111000) && ({row_reg, col_reg}<14'b11111010111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11111010111011) && ({row_reg, col_reg}<14'b11111010111101)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b11111010111101) && ({row_reg, col_reg}<14'b11111100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b11111100000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11111100000010) && ({row_reg, col_reg}<14'b11111100010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11111100010011) && ({row_reg, col_reg}<14'b11111100010110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11111100010110) && ({row_reg, col_reg}<14'b11111100011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b11111100011101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11111100011110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b11111100011111) && ({row_reg, col_reg}<14'b11111100100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b11111100100011) && ({row_reg, col_reg}<14'b11111100100101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b11111100100101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11111100100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b11111100100111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11111100101000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11111100101001) && ({row_reg, col_reg}<14'b11111100101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b11111100101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b11111100101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b11111100101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b11111100110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11111100110001) && ({row_reg, col_reg}<14'b11111100111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11111100111000) && ({row_reg, col_reg}<14'b11111100111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11111100111010) && ({row_reg, col_reg}<14'b11111100111101)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b11111100111101) && ({row_reg, col_reg}<14'b11111110000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b11111110000000) && ({row_reg, col_reg}<14'b11111110000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11111110000010) && ({row_reg, col_reg}<14'b11111110010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11111110010010) && ({row_reg, col_reg}<14'b11111110010110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11111110010110) && ({row_reg, col_reg}<14'b11111110011100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11111110011100) && ({row_reg, col_reg}<14'b11111110100001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b11111110100001) && ({row_reg, col_reg}<14'b11111110100101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b11111110100101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b11111110100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b11111110100111) && ({row_reg, col_reg}<14'b11111110101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b11111110101001) && ({row_reg, col_reg}<14'b11111110101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11111110101101) && ({row_reg, col_reg}<14'b11111110110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b11111110110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b11111110110001) && ({row_reg, col_reg}<14'b11111110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b11111110111000) && ({row_reg, col_reg}<14'b11111110111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b11111110111010) && ({row_reg, col_reg}<14'b11111110111101)) color_data = 12'b000100000000;

		if(({row_reg, col_reg}>=14'b11111110111101) && ({row_reg, col_reg}<=14'b11111111010111)) color_data = 12'b000000000000;
	end
endmodule