module shoot1_rom
	(
		input wire clk,
		input wire [5:0] row,
		input wire [6:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [5:0] row_reg;
	reg [6:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin
		if(({row_reg, col_reg}>=13'b0000000000000) && ({row_reg, col_reg}<13'b0000000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0000000100101) && ({row_reg, col_reg}<13'b0000000100111)) color_data = 12'b100000000000;

		if(({row_reg, col_reg}>=13'b0000000100111) && ({row_reg, col_reg}<13'b0000010100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0000010100100)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}>=13'b0000010100101) && ({row_reg, col_reg}<13'b0000010100111)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==13'b0000010100111)) color_data = 12'b011100000000;

		if(({row_reg, col_reg}>=13'b0000010101000) && ({row_reg, col_reg}<13'b0000100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0000100100011)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0000100100100)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}>=13'b0000100100101) && ({row_reg, col_reg}<13'b0000100100111)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0000100100111)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0000100101000)) color_data = 12'b011100000000;

		if(({row_reg, col_reg}>=13'b0000100101001) && ({row_reg, col_reg}<13'b0000110100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0000110100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0000110100010)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0000110100011)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0000110100100)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}>=13'b0000110100101) && ({row_reg, col_reg}<13'b0000110100111)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}==13'b0000110100111)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==13'b0000110101000)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0000110101001)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0000110101010)) color_data = 12'b001100110011;

		if(({row_reg, col_reg}>=13'b0000110101011) && ({row_reg, col_reg}<13'b0001000100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0001000100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001000100001)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0001000100010)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0001000100011)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==13'b0001000100100)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}>=13'b0001000100101) && ({row_reg, col_reg}<13'b0001000100111)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0001000100111)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0001000101000)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==13'b0001000101001)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0001000101010)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0001000101011)) color_data = 12'b001100110011;

		if(({row_reg, col_reg}>=13'b0001000101100) && ({row_reg, col_reg}<13'b0001010011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0001010011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0001010100000)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0001010100001)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0001010100010)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0001010100011)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==13'b0001010100100)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}>=13'b0001010100101) && ({row_reg, col_reg}<13'b0001010100111)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0001010100111)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}==13'b0001010101000)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==13'b0001010101001)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0001010101010)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0001010101011)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0001010101100)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=13'b0001010101101) && ({row_reg, col_reg}<13'b0001100011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0001100011111)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0001100100000)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0001100100001)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0001100100010)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0001100100011)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}==13'b0001100100100)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}>=13'b0001100100101) && ({row_reg, col_reg}<13'b0001100100111)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0001100100111)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0001100101000)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}==13'b0001100101001)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0001100101010)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0001100101011)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0001100101100)) color_data = 12'b011100000000;

		if(({row_reg, col_reg}>=13'b0001100101101) && ({row_reg, col_reg}<13'b0001110011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0001110011110)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0001110011111)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0001110100000)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0001110100001)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0001110100010)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}>=13'b0001110100011) && ({row_reg, col_reg}<13'b0001110101001)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0001110101001)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}==13'b0001110101010)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0001110101011)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0001110101100)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0001110101101)) color_data = 12'b011100000000;

		if(({row_reg, col_reg}>=13'b0001110101110) && ({row_reg, col_reg}<13'b0010000011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0010000011100)) color_data = 12'b011000000000;
		if(({row_reg, col_reg}==13'b0010000011101)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0010000011110)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0010000011111)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0010000100000)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}>=13'b0010000100001) && ({row_reg, col_reg}<13'b0010000100100)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0010000100100)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}>=13'b0010000100101) && ({row_reg, col_reg}<13'b0010000100111)) color_data = 12'b111100010001;
		if(({row_reg, col_reg}==13'b0010000100111)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}>=13'b0010000101000) && ({row_reg, col_reg}<13'b0010000101011)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0010000101011)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}==13'b0010000101100)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0010000101101)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0010000101110)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0010000101111)) color_data = 12'b011000000000;

		if(({row_reg, col_reg}>=13'b0010000110000) && ({row_reg, col_reg}<13'b0010010011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0010010011011) && ({row_reg, col_reg}<13'b0010010011101)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0010010011101)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0010010011110)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}>=13'b0010010011111) && ({row_reg, col_reg}<13'b0010010100010)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}==13'b0010010100010)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0010010100011)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0010010100100)) color_data = 12'b111100010001;
		if(({row_reg, col_reg}>=13'b0010010100101) && ({row_reg, col_reg}<13'b0010010100111)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}==13'b0010010100111)) color_data = 12'b111100010001;
		if(({row_reg, col_reg}==13'b0010010101000)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0010010101001)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}>=13'b0010010101010) && ({row_reg, col_reg}<13'b0010010101101)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}==13'b0010010101101)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==13'b0010010101110)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}>=13'b0010010101111) && ({row_reg, col_reg}<13'b0010010110001)) color_data = 12'b011100000000;

		if(({row_reg, col_reg}>=13'b0010010110001) && ({row_reg, col_reg}<13'b0010100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0010100011010) && ({row_reg, col_reg}<13'b0010100011100)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0010100011100)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0010100011101)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==13'b0010100011110)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0010100011111)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}==13'b0010100100000)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0010100100001)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}==13'b0010100100010)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0010100100011)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0010100100100)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}>=13'b0010100100101) && ({row_reg, col_reg}<13'b0010100100111)) color_data = 12'b111110011001;
		if(({row_reg, col_reg}==13'b0010100100111)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}==13'b0010100101000)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0010100101001)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0010100101010)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}==13'b0010100101011)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0010100101100)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}==13'b0010100101101)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0010100101110)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==13'b0010100101111)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}>=13'b0010100110000) && ({row_reg, col_reg}<13'b0010100110010)) color_data = 12'b011100000000;

		if(({row_reg, col_reg}>=13'b0010100110010) && ({row_reg, col_reg}<13'b0010110011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0010110011001)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0010110011010)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0010110011011)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==13'b0010110011100)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0010110011101)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}>=13'b0010110011110) && ({row_reg, col_reg}<13'b0010110100000)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}>=13'b0010110100000) && ({row_reg, col_reg}<13'b0010110100010)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0010110100010)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0010110100011)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}==13'b0010110100100)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}>=13'b0010110100101) && ({row_reg, col_reg}<13'b0010110100111)) color_data = 12'b111110111011;
		if(({row_reg, col_reg}==13'b0010110100111)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}==13'b0010110101000)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}==13'b0010110101001)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}>=13'b0010110101010) && ({row_reg, col_reg}<13'b0010110101100)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}>=13'b0010110101100) && ({row_reg, col_reg}<13'b0010110101110)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}==13'b0010110101110)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}==13'b0010110101111)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0010110110000)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==13'b0010110110001)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0010110110010)) color_data = 12'b011100000000;

		if(({row_reg, col_reg}>=13'b0010110110011) && ({row_reg, col_reg}<13'b0011000010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0011000010110)) color_data = 12'b011000000000;
		if(({row_reg, col_reg}>=13'b0011000010111) && ({row_reg, col_reg}<13'b0011000011001)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0011000011001)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0011000011010)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0011000011011)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}==13'b0011000011100)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}==13'b0011000011101)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0011000011110)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}==13'b0011000011111)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}>=13'b0011000100000) && ({row_reg, col_reg}<13'b0011000100010)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0011000100010)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}==13'b0011000100011)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}==13'b0011000100100)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}>=13'b0011000100101) && ({row_reg, col_reg}<13'b0011000100111)) color_data = 12'b111111011101;
		if(({row_reg, col_reg}==13'b0011000100111)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}==13'b0011000101000)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}==13'b0011000101001)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}>=13'b0011000101010) && ({row_reg, col_reg}<13'b0011000101100)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0011000101100)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0011000101101)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}==13'b0011000101110)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0011000101111)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}==13'b0011000110000)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}==13'b0011000110001)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0011000110010)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}>=13'b0011000110011) && ({row_reg, col_reg}<13'b0011000110101)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0011000110101)) color_data = 12'b011000000000;

		if(({row_reg, col_reg}>=13'b0011000110110) && ({row_reg, col_reg}<13'b0011010010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0011010010101)) color_data = 12'b011000000000;
		if(({row_reg, col_reg}==13'b0011010010110)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0011010010111)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0011010011000)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0011010011001)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0011010011010)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}>=13'b0011010011011) && ({row_reg, col_reg}<13'b0011010011110)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0011010011110)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}>=13'b0011010011111) && ({row_reg, col_reg}<13'b0011010100001)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0011010100001)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}==13'b0011010100010)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}==13'b0011010100011)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}==13'b0011010100100)) color_data = 12'b111110011001;
		if(({row_reg, col_reg}>=13'b0011010100101) && ({row_reg, col_reg}<13'b0011010100111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0011010100111)) color_data = 12'b111110011001;
		if(({row_reg, col_reg}==13'b0011010101000)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}==13'b0011010101001)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}==13'b0011010101010)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}>=13'b0011010101011) && ({row_reg, col_reg}<13'b0011010101101)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0011010101101)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}>=13'b0011010101110) && ({row_reg, col_reg}<13'b0011010110001)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0011010110001)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}==13'b0011010110010)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0011010110011)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0011010110100)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0011010110101)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0011010110110)) color_data = 12'b011000000000;

		if(({row_reg, col_reg}>=13'b0011010110111) && ({row_reg, col_reg}<13'b0011100010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0011100010101)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0011100010110)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0011100010111)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0011100011000)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}>=13'b0011100011001) && ({row_reg, col_reg}<13'b0011100011011)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}>=13'b0011100011011) && ({row_reg, col_reg}<13'b0011100011110)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0011100011110)) color_data = 12'b111100010001;
		if(({row_reg, col_reg}>=13'b0011100011111) && ({row_reg, col_reg}<13'b0011100100001)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}==13'b0011100100001)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}==13'b0011100100010)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}==13'b0011100100011)) color_data = 12'b111110011001;
		if(({row_reg, col_reg}==13'b0011100100100)) color_data = 12'b111111011100;
		if(({row_reg, col_reg}>=13'b0011100100101) && ({row_reg, col_reg}<13'b0011100100111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0011100100111)) color_data = 12'b111111011100;
		if(({row_reg, col_reg}==13'b0011100101000)) color_data = 12'b111110011001;
		if(({row_reg, col_reg}==13'b0011100101001)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}==13'b0011100101010)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}>=13'b0011100101011) && ({row_reg, col_reg}<13'b0011100101101)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}==13'b0011100101101)) color_data = 12'b111100010001;
		if(({row_reg, col_reg}>=13'b0011100101110) && ({row_reg, col_reg}<13'b0011100110001)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}>=13'b0011100110001) && ({row_reg, col_reg}<13'b0011100110011)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0011100110011)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}==13'b0011100110100)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0011100110101)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0011100110110)) color_data = 12'b011100000000;

		if(({row_reg, col_reg}>=13'b0011100110111) && ({row_reg, col_reg}<13'b0011110010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0011110010101)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0011110010110)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0011110010111)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}>=13'b0011110011000) && ({row_reg, col_reg}<13'b0011110011100)) color_data = 12'b111100010001;
		if(({row_reg, col_reg}>=13'b0011110011100) && ({row_reg, col_reg}<13'b0011110011111)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}>=13'b0011110011111) && ({row_reg, col_reg}<13'b0011110100001)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}==13'b0011110100001)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}==13'b0011110100010)) color_data = 12'b111110011001;
		if(({row_reg, col_reg}==13'b0011110100011)) color_data = 12'b111110111011;
		if(({row_reg, col_reg}==13'b0011110100100)) color_data = 12'b111111101101;
		if(({row_reg, col_reg}>=13'b0011110100101) && ({row_reg, col_reg}<13'b0011110100111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0011110100111)) color_data = 12'b111111101101;
		if(({row_reg, col_reg}==13'b0011110101000)) color_data = 12'b111110111011;
		if(({row_reg, col_reg}==13'b0011110101001)) color_data = 12'b111110011001;
		if(({row_reg, col_reg}==13'b0011110101010)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}>=13'b0011110101011) && ({row_reg, col_reg}<13'b0011110101101)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}>=13'b0011110101101) && ({row_reg, col_reg}<13'b0011110110000)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}>=13'b0011110110000) && ({row_reg, col_reg}<13'b0011110110100)) color_data = 12'b111100010001;
		if(({row_reg, col_reg}==13'b0011110110100)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==13'b0011110110101)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0011110110110)) color_data = 12'b011100000000;

		if(({row_reg, col_reg}>=13'b0011110110111) && ({row_reg, col_reg}<13'b0100000010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0100000010100)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0100000010101)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0100000010110)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0100000010111)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==13'b0100000011000)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0100000011001)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}>=13'b0100000011010) && ({row_reg, col_reg}<13'b0100000011100)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}>=13'b0100000011100) && ({row_reg, col_reg}<13'b0100000011111)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}>=13'b0100000011111) && ({row_reg, col_reg}<13'b0100000100001)) color_data = 12'b111110011001;
		if(({row_reg, col_reg}==13'b0100000100001)) color_data = 12'b111110111011;
		if(({row_reg, col_reg}==13'b0100000100010)) color_data = 12'b111111011100;
		if(({row_reg, col_reg}==13'b0100000100011)) color_data = 12'b111111011101;
		if(({row_reg, col_reg}>=13'b0100000100100) && ({row_reg, col_reg}<13'b0100000101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0100000101000)) color_data = 12'b111111011101;
		if(({row_reg, col_reg}==13'b0100000101001)) color_data = 12'b111111011100;
		if(({row_reg, col_reg}==13'b0100000101010)) color_data = 12'b111110111011;
		if(({row_reg, col_reg}>=13'b0100000101011) && ({row_reg, col_reg}<13'b0100000101101)) color_data = 12'b111110011001;
		if(({row_reg, col_reg}>=13'b0100000101101) && ({row_reg, col_reg}<13'b0100000110000)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}>=13'b0100000110000) && ({row_reg, col_reg}<13'b0100000110010)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}==13'b0100000110010)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}==13'b0100000110011)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0100000110100)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==13'b0100000110101)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0100000110110)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0100000110111)) color_data = 12'b011100000000;

		if(({row_reg, col_reg}>=13'b0100000111000) && ({row_reg, col_reg}<13'b0100010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0100010010100)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0100010010101)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0100010010110)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0100010010111)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0100010011000)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0100010011001)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}==13'b0100010011010)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}==13'b0100010011011)) color_data = 12'b111110101010;
		if(({row_reg, col_reg}==13'b0100010011100)) color_data = 12'b111110111011;
		if(({row_reg, col_reg}>=13'b0100010011101) && ({row_reg, col_reg}<13'b0100010011111)) color_data = 12'b111110101010;
		if(({row_reg, col_reg}==13'b0100010011111)) color_data = 12'b111110111011;
		if(({row_reg, col_reg}==13'b0100010100000)) color_data = 12'b111111011011;
		if(({row_reg, col_reg}==13'b0100010100001)) color_data = 12'b111111011101;
		if(({row_reg, col_reg}==13'b0100010100010)) color_data = 12'b111111101101;
		if(({row_reg, col_reg}>=13'b0100010100011) && ({row_reg, col_reg}<13'b0100010100101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=13'b0100010100101) && ({row_reg, col_reg}<13'b0100010100111)) color_data = 12'b111110111011;
		if(({row_reg, col_reg}>=13'b0100010100111) && ({row_reg, col_reg}<13'b0100010101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0100010101001)) color_data = 12'b111111101101;
		if(({row_reg, col_reg}==13'b0100010101010)) color_data = 12'b111111011101;
		if(({row_reg, col_reg}==13'b0100010101011)) color_data = 12'b111111011011;
		if(({row_reg, col_reg}==13'b0100010101100)) color_data = 12'b111110111011;
		if(({row_reg, col_reg}>=13'b0100010101101) && ({row_reg, col_reg}<13'b0100010101111)) color_data = 12'b111110101010;
		if(({row_reg, col_reg}==13'b0100010101111)) color_data = 12'b111110111011;
		if(({row_reg, col_reg}==13'b0100010110000)) color_data = 12'b111110101010;
		if(({row_reg, col_reg}==13'b0100010110001)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}==13'b0100010110010)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}==13'b0100010110011)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0100010110100)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0100010110101)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0100010110110)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0100010110111)) color_data = 12'b011100000000;

		if(({row_reg, col_reg}>=13'b0100010111000) && ({row_reg, col_reg}<13'b0100100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0100100010011) && ({row_reg, col_reg}<13'b0100100010101)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0100100010101)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0100100010110)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0100100010111)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}==13'b0100100011000)) color_data = 12'b111100010001;
		if(({row_reg, col_reg}==13'b0100100011001)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}==13'b0100100011010)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}==13'b0100100011011)) color_data = 12'b111110011001;
		if(({row_reg, col_reg}>=13'b0100100011100) && ({row_reg, col_reg}<13'b0100100011111)) color_data = 12'b111110111011;
		if(({row_reg, col_reg}==13'b0100100011111)) color_data = 12'b111111011100;
		if(({row_reg, col_reg}==13'b0100100100000)) color_data = 12'b111111011101;
		if(({row_reg, col_reg}==13'b0100100100001)) color_data = 12'b111111101101;
		if(({row_reg, col_reg}==13'b0100100100010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0100100100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0100100100100) && ({row_reg, col_reg}<13'b0100100100111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0100100100111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0100100101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0100100101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==13'b0100100101010)) color_data = 12'b111111101101;
		if(({row_reg, col_reg}==13'b0100100101011)) color_data = 12'b111111011101;
		if(({row_reg, col_reg}==13'b0100100101100)) color_data = 12'b111111011100;
		if(({row_reg, col_reg}>=13'b0100100101101) && ({row_reg, col_reg}<13'b0100100110000)) color_data = 12'b111110111011;
		if(({row_reg, col_reg}==13'b0100100110000)) color_data = 12'b111110011001;
		if(({row_reg, col_reg}==13'b0100100110001)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}==13'b0100100110010)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}==13'b0100100110011)) color_data = 12'b111100010001;
		if(({row_reg, col_reg}==13'b0100100110100)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}==13'b0100100110101)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0100100110110)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}>=13'b0100100110111) && ({row_reg, col_reg}<13'b0100100111001)) color_data = 12'b011100000000;

		if(({row_reg, col_reg}>=13'b0100100111001) && ({row_reg, col_reg}<13'b0100110010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0100110010011)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}>=13'b0100110010100) && ({row_reg, col_reg}<13'b0100110010110)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0100110010110)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0100110010111)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}==13'b0100110011000)) color_data = 12'b111100010001;
		if(({row_reg, col_reg}==13'b0100110011001)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}==13'b0100110011010)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}==13'b0100110011011)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}==13'b0100110011100)) color_data = 12'b111110101010;
		if(({row_reg, col_reg}==13'b0100110011101)) color_data = 12'b111110111011;
		if(({row_reg, col_reg}==13'b0100110011110)) color_data = 12'b111111011101;
		if(({row_reg, col_reg}>=13'b0100110011111) && ({row_reg, col_reg}<13'b0100110100001)) color_data = 12'b111111101101;
		if(({row_reg, col_reg}>=13'b0100110100001) && ({row_reg, col_reg}<13'b0100110100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0100110100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0100110100100) && ({row_reg, col_reg}<13'b0100110100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0100110100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b0100110100111) && ({row_reg, col_reg}<13'b0100110101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0100110101011) && ({row_reg, col_reg}<13'b0100110101101)) color_data = 12'b111111101101;
		if(({row_reg, col_reg}==13'b0100110101101)) color_data = 12'b111111011101;
		if(({row_reg, col_reg}==13'b0100110101110)) color_data = 12'b111110111011;
		if(({row_reg, col_reg}==13'b0100110101111)) color_data = 12'b111110101010;
		if(({row_reg, col_reg}==13'b0100110110000)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}==13'b0100110110001)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}==13'b0100110110010)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}==13'b0100110110011)) color_data = 12'b111100010001;
		if(({row_reg, col_reg}==13'b0100110110100)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}==13'b0100110110101)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}>=13'b0100110110110) && ({row_reg, col_reg}<13'b0100110111000)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0100110111000)) color_data = 12'b011100000000;

		if(({row_reg, col_reg}>=13'b0100110111001) && ({row_reg, col_reg}<13'b0101000010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0101000010010) && ({row_reg, col_reg}<13'b0101000010100)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}>=13'b0101000010100) && ({row_reg, col_reg}<13'b0101000010111)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0101000010111)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}>=13'b0101000011000) && ({row_reg, col_reg}<13'b0101000011010)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}==13'b0101000011010)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}==13'b0101000011011)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}==13'b0101000011100)) color_data = 12'b111110101010;
		if(({row_reg, col_reg}==13'b0101000011101)) color_data = 12'b111111011011;
		if(({row_reg, col_reg}==13'b0101000011110)) color_data = 12'b111111101101;
		if(({row_reg, col_reg}>=13'b0101000011111) && ({row_reg, col_reg}<13'b0101000100001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=13'b0101000100001) && ({row_reg, col_reg}<13'b0101000100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0101000100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0101000100100) && ({row_reg, col_reg}<13'b0101000100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0101000100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b0101000100111) && ({row_reg, col_reg}<13'b0101000101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0101000101001) && ({row_reg, col_reg}<13'b0101000101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0101000101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0101000101100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0101000101101)) color_data = 12'b111111101101;
		if(({row_reg, col_reg}==13'b0101000101110)) color_data = 12'b111111011011;
		if(({row_reg, col_reg}==13'b0101000101111)) color_data = 12'b111110101010;
		if(({row_reg, col_reg}==13'b0101000110000)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}==13'b0101000110001)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}>=13'b0101000110010) && ({row_reg, col_reg}<13'b0101000110100)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}==13'b0101000110100)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}>=13'b0101000110101) && ({row_reg, col_reg}<13'b0101000111000)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}>=13'b0101000111000) && ({row_reg, col_reg}<13'b0101000111010)) color_data = 12'b011100000000;

		if(({row_reg, col_reg}>=13'b0101000111010) && ({row_reg, col_reg}<13'b0101010010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0101010010001) && ({row_reg, col_reg}<13'b0101010010011)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0101010010011)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}>=13'b0101010010100) && ({row_reg, col_reg}<13'b0101010010110)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0101010010110)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==13'b0101010010111)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0101010011000)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}==13'b0101010011001)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}==13'b0101010011010)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}==13'b0101010011011)) color_data = 12'b111110011001;
		if(({row_reg, col_reg}==13'b0101010011100)) color_data = 12'b111110111011;
		if(({row_reg, col_reg}==13'b0101010011101)) color_data = 12'b111111011101;
		if(({row_reg, col_reg}>=13'b0101010011110) && ({row_reg, col_reg}<13'b0101010100000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==13'b0101010100000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0101010100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0101010100010) && ({row_reg, col_reg}<13'b0101010100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0101010100100) && ({row_reg, col_reg}<13'b0101010100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0101010100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0101010100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0101010101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0101010101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=13'b0101010101010) && ({row_reg, col_reg}<13'b0101010101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0101010101100) && ({row_reg, col_reg}<13'b0101010101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0101010101110)) color_data = 12'b111111011101;
		if(({row_reg, col_reg}==13'b0101010101111)) color_data = 12'b111110111011;
		if(({row_reg, col_reg}==13'b0101010110000)) color_data = 12'b111110011001;
		if(({row_reg, col_reg}==13'b0101010110001)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}==13'b0101010110010)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}==13'b0101010110011)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}==13'b0101010110100)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0101010110101)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}>=13'b0101010110110) && ({row_reg, col_reg}<13'b0101010111000)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0101010111000)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}>=13'b0101010111001) && ({row_reg, col_reg}<13'b0101010111011)) color_data = 12'b011100000000;

		if(({row_reg, col_reg}>=13'b0101010111011) && ({row_reg, col_reg}<13'b0101100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0101100010000)) color_data = 12'b011000000000;
		if(({row_reg, col_reg}>=13'b0101100010001) && ({row_reg, col_reg}<13'b0101100010011)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}>=13'b0101100010011) && ({row_reg, col_reg}<13'b0101100010110)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==13'b0101100010110)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0101100010111)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0101100011000)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0101100011001)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}==13'b0101100011010)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}==13'b0101100011011)) color_data = 12'b111110101010;
		if(({row_reg, col_reg}==13'b0101100011100)) color_data = 12'b111111011101;
		if(({row_reg, col_reg}>=13'b0101100011101) && ({row_reg, col_reg}<13'b0101100011111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==13'b0101100011111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=13'b0101100100000) && ({row_reg, col_reg}<13'b0101100100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0101100100010) && ({row_reg, col_reg}<13'b0101100100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0101100100100) && ({row_reg, col_reg}<13'b0101100100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0101100100110) && ({row_reg, col_reg}<13'b0101100101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0101100101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0101100101001) && ({row_reg, col_reg}<13'b0101100101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0101100101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0101100101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0101100101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0101100101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0101100101111)) color_data = 12'b111111011101;
		if(({row_reg, col_reg}==13'b0101100110000)) color_data = 12'b111110101010;
		if(({row_reg, col_reg}==13'b0101100110001)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}==13'b0101100110010)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}==13'b0101100110011)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0101100110100)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0101100110101)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}>=13'b0101100110110) && ({row_reg, col_reg}<13'b0101100111001)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}>=13'b0101100111001) && ({row_reg, col_reg}<13'b0101100111011)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0101100111011)) color_data = 12'b011000000000;

		if(({row_reg, col_reg}>=13'b0101100111100) && ({row_reg, col_reg}<13'b0101110001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0101110001111)) color_data = 12'b011000000000;
		if(({row_reg, col_reg}>=13'b0101110010000) && ({row_reg, col_reg}<13'b0101110010010)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0101110010010)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}>=13'b0101110010011) && ({row_reg, col_reg}<13'b0101110010101)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0101110010101)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}==13'b0101110010110)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}>=13'b0101110010111) && ({row_reg, col_reg}<13'b0101110011001)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0101110011001)) color_data = 12'b111100010001;
		if(({row_reg, col_reg}==13'b0101110011010)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}==13'b0101110011011)) color_data = 12'b111110111011;
		if(({row_reg, col_reg}==13'b0101110011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=13'b0101110011101) && ({row_reg, col_reg}<13'b0101110100000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=13'b0101110100000) && ({row_reg, col_reg}<13'b0101110100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0101110100010) && ({row_reg, col_reg}<13'b0101110100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0101110100100) && ({row_reg, col_reg}<13'b0101110100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0101110100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0101110100111) && ({row_reg, col_reg}<13'b0101110101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0101110101001) && ({row_reg, col_reg}<13'b0101110101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0101110101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0101110101100) && ({row_reg, col_reg}<13'b0101110101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0101110101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0101110101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0101110110000)) color_data = 12'b111110111011;
		if(({row_reg, col_reg}==13'b0101110110001)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}==13'b0101110110010)) color_data = 12'b111100010001;
		if(({row_reg, col_reg}>=13'b0101110110011) && ({row_reg, col_reg}<13'b0101110110101)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0101110110101)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0101110110110)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}>=13'b0101110110111) && ({row_reg, col_reg}<13'b0101110111001)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0101110111001)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}>=13'b0101110111010) && ({row_reg, col_reg}<13'b0101110111100)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0101110111100)) color_data = 12'b011000000000;

		if(({row_reg, col_reg}>=13'b0101110111101) && ({row_reg, col_reg}<13'b0110000001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0110000001110)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0110000001111)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0110000010000)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==13'b0110000010001)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0110000010010)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}>=13'b0110000010011) && ({row_reg, col_reg}<13'b0110000010101)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}==13'b0110000010101)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0110000010110)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}>=13'b0110000010111) && ({row_reg, col_reg}<13'b0110000011001)) color_data = 12'b111100010001;
		if(({row_reg, col_reg}==13'b0110000011001)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}==13'b0110000011010)) color_data = 12'b111110011001;
		if(({row_reg, col_reg}==13'b0110000011011)) color_data = 12'b111111011100;
		if(({row_reg, col_reg}==13'b0110000011100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=13'b0110000011101) && ({row_reg, col_reg}<13'b0110000011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0110000011111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=13'b0110000100000) && ({row_reg, col_reg}<13'b0110000100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0110000100010) && ({row_reg, col_reg}<13'b0110000100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0110000100100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0110000100101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0110000100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b0110000100111) && ({row_reg, col_reg}<13'b0110000101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0110000101001) && ({row_reg, col_reg}<13'b0110000101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0110000101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0110000101100) && ({row_reg, col_reg}<13'b0110000101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0110000101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0110000110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110000110001)) color_data = 12'b111110011001;
		if(({row_reg, col_reg}==13'b0110000110010)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}>=13'b0110000110011) && ({row_reg, col_reg}<13'b0110000110101)) color_data = 12'b111100010001;
		if(({row_reg, col_reg}==13'b0110000110101)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0110000110110)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}>=13'b0110000110111) && ({row_reg, col_reg}<13'b0110000111001)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}==13'b0110000111001)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}==13'b0110000111010)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0110000111011)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==13'b0110000111100)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0110000111101)) color_data = 12'b011100000000;

		if(({row_reg, col_reg}>=13'b0110000111110) && ({row_reg, col_reg}<13'b0110010001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0110010001100)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0110010001101)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0110010001110)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}>=13'b0110010001111) && ({row_reg, col_reg}<13'b0110010010001)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0110010010001)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}>=13'b0110010010010) && ({row_reg, col_reg}<13'b0110010010100)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}>=13'b0110010010100) && ({row_reg, col_reg}<13'b0110010010111)) color_data = 12'b111100010001;
		if(({row_reg, col_reg}==13'b0110010010111)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}==13'b0110010011000)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}==13'b0110010011001)) color_data = 12'b111110011001;
		if(({row_reg, col_reg}==13'b0110010011010)) color_data = 12'b111110111011;
		if(({row_reg, col_reg}>=13'b0110010011011) && ({row_reg, col_reg}<13'b0110010011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0110010011101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==13'b0110010011110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==13'b0110010011111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=13'b0110010100000) && ({row_reg, col_reg}<13'b0110010100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0110010100010) && ({row_reg, col_reg}<13'b0110010100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0110010100100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0110010100101) && ({row_reg, col_reg}<13'b0110010100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0110010100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0110010101000) && ({row_reg, col_reg}<13'b0110010101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0110010101100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0110010101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0110010101110) && ({row_reg, col_reg}<13'b0110010110000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b0110010110000) && ({row_reg, col_reg}<13'b0110010110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110010110010)) color_data = 12'b111110011001;
		if(({row_reg, col_reg}==13'b0110010110011)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}==13'b0110010110100)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}>=13'b0110010110101) && ({row_reg, col_reg}<13'b0110010111000)) color_data = 12'b111100010001;
		if(({row_reg, col_reg}>=13'b0110010111000) && ({row_reg, col_reg}<13'b0110010111010)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0110010111010)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}>=13'b0110010111011) && ({row_reg, col_reg}<13'b0110010111101)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0110010111101)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0110010111110)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0110010111111)) color_data = 12'b011100000000;

		if(({row_reg, col_reg}>=13'b0110011000000) && ({row_reg, col_reg}<13'b0110100001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0110100001001)) color_data = 12'b011000000000;
		if(({row_reg, col_reg}>=13'b0110100001010) && ({row_reg, col_reg}<13'b0110100001100)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0110100001100)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==13'b0110100001101)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}>=13'b0110100001110) && ({row_reg, col_reg}<13'b0110100010001)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0110100010001)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}>=13'b0110100010010) && ({row_reg, col_reg}<13'b0110100010101)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}>=13'b0110100010101) && ({row_reg, col_reg}<13'b0110100010111)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}==13'b0110100010111)) color_data = 12'b111110011001;
		if(({row_reg, col_reg}==13'b0110100011000)) color_data = 12'b111110101010;
		if(({row_reg, col_reg}==13'b0110100011001)) color_data = 12'b111111011011;
		if(({row_reg, col_reg}>=13'b0110100011010) && ({row_reg, col_reg}<13'b0110100011100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==13'b0110100011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=13'b0110100011101) && ({row_reg, col_reg}<13'b0110100011111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=13'b0110100011111) && ({row_reg, col_reg}<13'b0110100100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0110100100010) && ({row_reg, col_reg}<13'b0110100100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0110100100100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0110100100101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0110100100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0110100100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0110100101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0110100101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=13'b0110100101010) && ({row_reg, col_reg}<13'b0110100101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0110100101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0110100101101) && ({row_reg, col_reg}<13'b0110100110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110100110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0110100110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110100110010)) color_data = 12'b111111011011;
		if(({row_reg, col_reg}==13'b0110100110011)) color_data = 12'b111110101010;
		if(({row_reg, col_reg}==13'b0110100110100)) color_data = 12'b111110011001;
		if(({row_reg, col_reg}>=13'b0110100110101) && ({row_reg, col_reg}<13'b0110100110111)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}>=13'b0110100110111) && ({row_reg, col_reg}<13'b0110100111010)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}==13'b0110100111010)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}>=13'b0110100111011) && ({row_reg, col_reg}<13'b0110100111110)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0110100111110)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}==13'b0110100111111)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}>=13'b0110101000000) && ({row_reg, col_reg}<13'b0110101000010)) color_data = 12'b011100000000;

		if(({row_reg, col_reg}==13'b0110101000010)) color_data = 12'b011000000000;
		if(({row_reg, col_reg}>=13'b0110110000000) && ({row_reg, col_reg}<13'b0110110001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0110110001001)) color_data = 12'b011000000000;
		if(({row_reg, col_reg}==13'b0110110001010)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0110110001011)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0110110001100)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==13'b0110110001101)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}==13'b0110110001110)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}>=13'b0110110001111) && ({row_reg, col_reg}<13'b0110110010001)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}>=13'b0110110010001) && ({row_reg, col_reg}<13'b0110110010100)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}>=13'b0110110010100) && ({row_reg, col_reg}<13'b0110110010111)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}==13'b0110110010111)) color_data = 12'b111110011001;
		if(({row_reg, col_reg}==13'b0110110011000)) color_data = 12'b111110111011;
		if(({row_reg, col_reg}==13'b0110110011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0110110011010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==13'b0110110011011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==13'b0110110011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=13'b0110110011101) && ({row_reg, col_reg}<13'b0110110011111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=13'b0110110011111) && ({row_reg, col_reg}<13'b0110110100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0110110100001) && ({row_reg, col_reg}<13'b0110110100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0110110100100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0110110100101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0110110100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0110110100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0110110101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0110110101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=13'b0110110101010) && ({row_reg, col_reg}<13'b0110110101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0110110101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0110110101101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0110110101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0110110101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0110110110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0110110110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0110110110011)) color_data = 12'b111110111011;
		if(({row_reg, col_reg}==13'b0110110110100)) color_data = 12'b111110011001;
		if(({row_reg, col_reg}>=13'b0110110110101) && ({row_reg, col_reg}<13'b0110110111000)) color_data = 12'b111101110111;
		if(({row_reg, col_reg}>=13'b0110110111000) && ({row_reg, col_reg}<13'b0110110111011)) color_data = 12'b111101010101;
		if(({row_reg, col_reg}>=13'b0110110111011) && ({row_reg, col_reg}<13'b0110110111101)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0110110111101)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}==13'b0110110111110)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}==13'b0110110111111)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==13'b0110111000000)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0110111000001)) color_data = 12'b011100000000;

		if(({row_reg, col_reg}==13'b0110111000010)) color_data = 12'b011000000000;
		if(({row_reg, col_reg}>=13'b0111000000000) && ({row_reg, col_reg}<13'b0111000001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0111000001100)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}>=13'b0111000001101) && ({row_reg, col_reg}<13'b0111000001111)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}>=13'b0111000001111) && ({row_reg, col_reg}<13'b0111000010001)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}>=13'b0111000010001) && ({row_reg, col_reg}<13'b0111000010011)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0111000010011)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}==13'b0111000010100)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0111000010101)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0111000010110)) color_data = 12'b111100010001;
		if(({row_reg, col_reg}==13'b0111000010111)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}==13'b0111000011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111000011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0111000011010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=13'b0111000011011) && ({row_reg, col_reg}<13'b0111000011101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==13'b0111000011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0111000011110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=13'b0111000011111) && ({row_reg, col_reg}<13'b0111000100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0111000100001) && ({row_reg, col_reg}<13'b0111000100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0111000100011) && ({row_reg, col_reg}<13'b0111000100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0111000100101) && ({row_reg, col_reg}<13'b0111000100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0111000100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0111000101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0111000101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0111000101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0111000101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0111000101100) && ({row_reg, col_reg}<13'b0111000101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0111000101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0111000101111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0111000110000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0111000110001) && ({row_reg, col_reg}<13'b0111000110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0111000110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111000110100)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}==13'b0111000110101)) color_data = 12'b111100010001;
		if(({row_reg, col_reg}==13'b0111000110110)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0111000110111)) color_data = 12'b111000000000;
		if(({row_reg, col_reg}==13'b0111000111000)) color_data = 12'b110100000000;
		if(({row_reg, col_reg}>=13'b0111000111001) && ({row_reg, col_reg}<13'b0111000111011)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}>=13'b0111000111011) && ({row_reg, col_reg}<13'b0111000111101)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}>=13'b0111000111101) && ({row_reg, col_reg}<13'b0111000111111)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0111000111111)) color_data = 12'b011100000000;

		if(({row_reg, col_reg}>=13'b0111001000000) && ({row_reg, col_reg}<13'b0111010001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0111010001111) && ({row_reg, col_reg}<13'b0111010010010)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}>=13'b0111010010010) && ({row_reg, col_reg}<13'b0111010010100)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0111010010100)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0111010010101)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}==13'b0111010010110)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0111010010111)) color_data = 12'b111100010001;
		if(({row_reg, col_reg}==13'b0111010011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111010011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b0111010011010) && ({row_reg, col_reg}<13'b0111010011100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=13'b0111010011100) && ({row_reg, col_reg}<13'b0111010011110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0111010011110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=13'b0111010011111) && ({row_reg, col_reg}<13'b0111010100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0111010100001) && ({row_reg, col_reg}<13'b0111010100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0111010100011) && ({row_reg, col_reg}<13'b0111010100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0111010100101) && ({row_reg, col_reg}<13'b0111010100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0111010100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=13'b0111010101000) && ({row_reg, col_reg}<13'b0111010101011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0111010101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0111010101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b0111010101101) && ({row_reg, col_reg}<13'b0111010110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0111010110000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0111010110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0111010110010) && ({row_reg, col_reg}<13'b0111010110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0111010110100)) color_data = 12'b111100010001;
		if(({row_reg, col_reg}==13'b0111010110101)) color_data = 12'b111100000000;
		if(({row_reg, col_reg}==13'b0111010110110)) color_data = 12'b110000000000;
		if(({row_reg, col_reg}==13'b0111010110111)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}>=13'b0111010111000) && ({row_reg, col_reg}<13'b0111010111010)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}>=13'b0111010111010) && ({row_reg, col_reg}<13'b0111010111101)) color_data = 12'b011100000000;

		if(({row_reg, col_reg}>=13'b0111010111101) && ({row_reg, col_reg}<13'b0111100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b0111100010001)) color_data = 12'b011000000000;
		if(({row_reg, col_reg}==13'b0111100010010)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}>=13'b0111100010011) && ({row_reg, col_reg}<13'b0111100010101)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0111100010101)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0111100010110)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0111100010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111100011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0111100011001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=13'b0111100011010) && ({row_reg, col_reg}<13'b0111100011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b0111100011100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==13'b0111100011101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==13'b0111100011110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=13'b0111100011111) && ({row_reg, col_reg}<13'b0111100100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0111100100001) && ({row_reg, col_reg}<13'b0111100100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b0111100100011) && ({row_reg, col_reg}<13'b0111100100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b0111100100101) && ({row_reg, col_reg}<13'b0111100100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0111100100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=13'b0111100101000) && ({row_reg, col_reg}<13'b0111100101011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0111100101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0111100101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0111100101101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b0111100101110) && ({row_reg, col_reg}<13'b0111100110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0111100110000) && ({row_reg, col_reg}<13'b0111100110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0111100110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0111100110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111100110101)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==13'b0111100110110)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}>=13'b0111100110111) && ({row_reg, col_reg}<13'b0111100111001)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0111100111001)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0111100111010)) color_data = 12'b011000000000;

		if(({row_reg, col_reg}>=13'b0111100111011) && ({row_reg, col_reg}<13'b0111110010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0111110010010) && ({row_reg, col_reg}<13'b0111110010100)) color_data = 12'b011000000000;
		if(({row_reg, col_reg}==13'b0111110010100)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b0111110010101)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0111110010110)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==13'b0111110010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111110011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b0111110011001) && ({row_reg, col_reg}<13'b0111110011011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==13'b0111110011011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=13'b0111110011100) && ({row_reg, col_reg}<13'b0111110011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0111110011110) && ({row_reg, col_reg}<13'b0111110100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b0111110100001) && ({row_reg, col_reg}<13'b0111110100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b0111110100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b0111110100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0111110100101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b0111110100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0111110100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=13'b0111110101000) && ({row_reg, col_reg}<13'b0111110101011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b0111110101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b0111110101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b0111110101101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b0111110101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111110101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b0111110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b0111110110001) && ({row_reg, col_reg}<13'b0111110110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111110110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b0111110110100) && ({row_reg, col_reg}<13'b0111110110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b0111110110110)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==13'b0111110110111)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}>=13'b0111110111000) && ({row_reg, col_reg}<13'b0111110111010)) color_data = 12'b011000000000;

		if(({row_reg, col_reg}>=13'b0111110111010) && ({row_reg, col_reg}<13'b1000000010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1000000010100)) color_data = 12'b011000000000;
		if(({row_reg, col_reg}==13'b1000000010101)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b1000000010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1000000010111) && ({row_reg, col_reg}<13'b1000000011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1000000011001) && ({row_reg, col_reg}<13'b1000000011011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=13'b1000000011011) && ({row_reg, col_reg}<13'b1000000011110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=13'b1000000011110) && ({row_reg, col_reg}<13'b1000000100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1000000100001) && ({row_reg, col_reg}<13'b1000000100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1000000100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1000000100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1000000100101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b1000000100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b1000000100111) && ({row_reg, col_reg}<13'b1000000101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=13'b1000000101001) && ({row_reg, col_reg}<13'b1000000101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b1000000101011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=13'b1000000101100) && ({row_reg, col_reg}<13'b1000000101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b1000000101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b1000000101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1000000110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1000000110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b1000000110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1000000110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1000000110100) && ({row_reg, col_reg}<13'b1000000110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1000000110110)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==13'b1000000110111)) color_data = 12'b011000000000;

		if(({row_reg, col_reg}>=13'b1000000111000) && ({row_reg, col_reg}<13'b1000010010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1000010010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b1000010010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1000010010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b1000010011000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==13'b1000010011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=13'b1000010011010) && ({row_reg, col_reg}<13'b1000010011100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b1000010011100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==13'b1000010011101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=13'b1000010011110) && ({row_reg, col_reg}<13'b1000010100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1000010100001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1000010100010) && ({row_reg, col_reg}<13'b1000010100100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1000010100100) && ({row_reg, col_reg}<13'b1000010100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b1000010100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b1000010100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=13'b1000010101000) && ({row_reg, col_reg}<13'b1000010101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b1000010101011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b1000010101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=13'b1000010101101) && ({row_reg, col_reg}<13'b1000010101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b1000010101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b1000010110000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1000010110001) && ({row_reg, col_reg}<13'b1000010110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1000010110011) && ({row_reg, col_reg}<13'b1000010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1000010110101) && ({row_reg, col_reg}<13'b1000010110111)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=13'b1000010110111) && ({row_reg, col_reg}<13'b1000100010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b1000100010101) && ({row_reg, col_reg}<13'b1000100010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1000100010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b1000100011000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=13'b1000100011001) && ({row_reg, col_reg}<13'b1000100011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b1000100011011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=13'b1000100011100) && ({row_reg, col_reg}<13'b1000100011110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=13'b1000100011110) && ({row_reg, col_reg}<13'b1000100100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1000100100001) && ({row_reg, col_reg}<13'b1000100100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1000100100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1000100100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b1000100100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b1000100100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b1000100100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=13'b1000100101000) && ({row_reg, col_reg}<13'b1000100101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b1000100101011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b1000100101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b1000100101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b1000100101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1000100101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1000100110000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1000100110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1000100110010) && ({row_reg, col_reg}<13'b1000100110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1000100110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1000100110101) && ({row_reg, col_reg}<13'b1000100110111)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=13'b1000100110111) && ({row_reg, col_reg}<13'b1000110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1000110010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1000110010101) && ({row_reg, col_reg}<13'b1000110010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1000110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b1000110011000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==13'b1000110011001)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==13'b1000110011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b1000110011011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=13'b1000110011100) && ({row_reg, col_reg}<13'b1000110011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b1000110011110) && ({row_reg, col_reg}<13'b1000110100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1000110100000) && ({row_reg, col_reg}<13'b1000110100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1000110100010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1000110100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1000110100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b1000110100101) && ({row_reg, col_reg}<13'b1000110100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b1000110100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b1000110101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=13'b1000110101001) && ({row_reg, col_reg}<13'b1000110101011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==13'b1000110101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b1000110101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b1000110101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b1000110101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1000110101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b1000110110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1000110110001) && ({row_reg, col_reg}<13'b1000110110011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1000110110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1000110110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1000110110101) && ({row_reg, col_reg}<13'b1000110111000)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=13'b1000110111000) && ({row_reg, col_reg}<13'b1001000010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b1001000010100) && ({row_reg, col_reg}<13'b1001000010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1001000010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b1001000010111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=13'b1001000011000) && ({row_reg, col_reg}<13'b1001000011010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b1001000011010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==13'b1001000011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1001000011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==13'b1001000011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1001000011110) && ({row_reg, col_reg}<13'b1001000100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1001000100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1001000100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1001000100010) && ({row_reg, col_reg}<13'b1001000100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1001000100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b1001000100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b1001000100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==13'b1001000100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=13'b1001000101000) && ({row_reg, col_reg}<13'b1001000101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==13'b1001000101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b1001000101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b1001000101110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1001000101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1001000110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1001000110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b1001000110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1001000110011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1001000110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1001000110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1001000110110) && ({row_reg, col_reg}<13'b1001000111000)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=13'b1001000111000) && ({row_reg, col_reg}<13'b1001010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1001010010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1001010010101) && ({row_reg, col_reg}<13'b1001010010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b1001010010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b1001010011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==13'b1001010011001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==13'b1001010011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1001010011011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==13'b1001010011100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=13'b1001010011101) && ({row_reg, col_reg}<13'b1001010100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1001010100001) && ({row_reg, col_reg}<13'b1001010100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1001010100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1001010100100) && ({row_reg, col_reg}<13'b1001010100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1001010100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b1001010100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=13'b1001010101000) && ({row_reg, col_reg}<13'b1001010101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==13'b1001010101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b1001010101101) && ({row_reg, col_reg}<13'b1001010110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b1001010110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1001010110001) && ({row_reg, col_reg}<13'b1001010110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b1001010110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1001010110101) && ({row_reg, col_reg}<13'b1001010110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b1001010110111)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=13'b1001010111000) && ({row_reg, col_reg}<13'b1001100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b1001100010011) && ({row_reg, col_reg}<13'b1001100010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1001100010101) && ({row_reg, col_reg}<13'b1001100101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1001100101111) && ({row_reg, col_reg}<13'b1001100110011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1001100110011) && ({row_reg, col_reg}<13'b1001100110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1001100110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b1001100111000)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=13'b1001100111001) && ({row_reg, col_reg}<13'b1001110010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b1001110010011) && ({row_reg, col_reg}<13'b1001110010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1001110010101) && ({row_reg, col_reg}<13'b1001110011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1001110011011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1001110011100) && ({row_reg, col_reg}<13'b1001110100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1001110100001) && ({row_reg, col_reg}<13'b1001110110011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1001110110011) && ({row_reg, col_reg}<13'b1001110110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1001110110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1001110110111) && ({row_reg, col_reg}<13'b1001110111001)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=13'b1001110111001) && ({row_reg, col_reg}<13'b1010000010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1010000010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1010000010100) && ({row_reg, col_reg}<13'b1010000100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1010000100001) && ({row_reg, col_reg}<13'b1010000101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1010000101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1010000110000) && ({row_reg, col_reg}<13'b1010000110011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1010000110011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1010000110100) && ({row_reg, col_reg}<13'b1010000110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1010000110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1010000110111) && ({row_reg, col_reg}<13'b1010000111001)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=13'b1010000111001) && ({row_reg, col_reg}<13'b1010010010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b1010010010010) && ({row_reg, col_reg}<13'b1010010010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1010010010100) && ({row_reg, col_reg}<13'b1010010100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1010010100001) && ({row_reg, col_reg}<13'b1010010101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1010010101111) && ({row_reg, col_reg}<13'b1010010110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1010010110001) && ({row_reg, col_reg}<13'b1010010110011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1010010110011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1010010110100) && ({row_reg, col_reg}<13'b1010010110111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1010010110111) && ({row_reg, col_reg}<13'b1010010111010)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=13'b1010010111010) && ({row_reg, col_reg}<13'b1010100010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1010100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1010100010011) && ({row_reg, col_reg}<13'b1010100011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1010100011101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1010100011110) && ({row_reg, col_reg}<13'b1010100100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1010100100001) && ({row_reg, col_reg}<13'b1010100101011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1010100101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1010100101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1010100101101) && ({row_reg, col_reg}<13'b1010100110000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1010100110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1010100110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1010100110010) && ({row_reg, col_reg}<13'b1010100110100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1010100110100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1010100110101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1010100110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1010100110111) && ({row_reg, col_reg}<13'b1010100111010)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=13'b1010100111010) && ({row_reg, col_reg}<13'b1010110010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1010110010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1010110010010) && ({row_reg, col_reg}<13'b1010110010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1010110010101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1010110010110) && ({row_reg, col_reg}<13'b1010110100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1010110100000) && ({row_reg, col_reg}<13'b1010110101011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1010110101011) && ({row_reg, col_reg}<13'b1010110110011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1010110110011) && ({row_reg, col_reg}<13'b1010110110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1010110110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1010110110111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1010110111000) && ({row_reg, col_reg}<13'b1010110111011)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=13'b1010110111011) && ({row_reg, col_reg}<13'b1011000010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1011000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1011000010010) && ({row_reg, col_reg}<13'b1011000010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1011000010101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1011000010110) && ({row_reg, col_reg}<13'b1011000011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1011000011111) && ({row_reg, col_reg}<13'b1011000101001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1011000101001) && ({row_reg, col_reg}<13'b1011000110011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1011000110011) && ({row_reg, col_reg}<13'b1011000110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1011000110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1011000110111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1011000111000) && ({row_reg, col_reg}<13'b1011000111011)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=13'b1011000111011) && ({row_reg, col_reg}<13'b1011010010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1011010010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1011010010001) && ({row_reg, col_reg}<13'b1011010010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1011010010100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1011010010101) && ({row_reg, col_reg}<13'b1011010011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1011010011100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1011010011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1011010011110) && ({row_reg, col_reg}<13'b1011010100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1011010100010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1011010100011) && ({row_reg, col_reg}<13'b1011010100111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1011010100111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1011010101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1011010101001) && ({row_reg, col_reg}<13'b1011010110100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1011010110100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1011010110101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1011010110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1011010110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1011010111000) && ({row_reg, col_reg}<13'b1011010111100)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=13'b1011010111100) && ({row_reg, col_reg}<13'b1011100001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b1011100001111) && ({row_reg, col_reg}<13'b1011100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1011100010001) && ({row_reg, col_reg}<13'b1011100011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1011100011100) && ({row_reg, col_reg}<13'b1011100100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1011100100010) && ({row_reg, col_reg}<13'b1011100110101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1011100110101) && ({row_reg, col_reg}<13'b1011100111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1011100111001) && ({row_reg, col_reg}<13'b1011100111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1011100111100)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=13'b1011100111101) && ({row_reg, col_reg}<13'b1011110001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b1011110001111) && ({row_reg, col_reg}<13'b1011110010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1011110010001) && ({row_reg, col_reg}<13'b1011110010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1011110010110) && ({row_reg, col_reg}<13'b1011110011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1011110011000) && ({row_reg, col_reg}<13'b1011110011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1011110011010) && ({row_reg, col_reg}<13'b1011110100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1011110100010) && ({row_reg, col_reg}<13'b1011110110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1011110110111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1011110111000) && ({row_reg, col_reg}<13'b1011110111101)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=13'b1011110111101) && ({row_reg, col_reg}<13'b1100000001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1100000001100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==13'b1100000001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b1100000001110) && ({row_reg, col_reg}<13'b1100000010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1100000010000) && ({row_reg, col_reg}<13'b1100000010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1100000010101) && ({row_reg, col_reg}<13'b1100000100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1100000100000) && ({row_reg, col_reg}<13'b1100000111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1100000111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1100000111001) && ({row_reg, col_reg}<13'b1100000111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1100000111101)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=13'b1100000111110) && ({row_reg, col_reg}<13'b1100010001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1100010001011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==13'b1100010001100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b1100010001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1100010001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1100010001111) && ({row_reg, col_reg}<13'b1100010010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1100010010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b1100010010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1100010010100) && ({row_reg, col_reg}<13'b1100010011110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1100010011110) && ({row_reg, col_reg}<13'b1100010110000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1100010110000) && ({row_reg, col_reg}<13'b1100010110010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b1100010110010) && ({row_reg, col_reg}<13'b1100010110100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1100010110100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b1100010110101) && ({row_reg, col_reg}<13'b1100010110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1100010110111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1100010111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1100010111001) && ({row_reg, col_reg}<13'b1100010111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1100010111101)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=13'b1100010111110) && ({row_reg, col_reg}<13'b1100100001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=13'b1100100001001) && ({row_reg, col_reg}<13'b1100100001011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==13'b1100100001011)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==13'b1100100001100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=13'b1100100001101) && ({row_reg, col_reg}<13'b1100100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b1100100010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1100100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1100100010010) && ({row_reg, col_reg}<13'b1100100010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1100100010110) && ({row_reg, col_reg}<13'b1100100011101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1100100011101) && ({row_reg, col_reg}<13'b1100100101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1100100101111) && ({row_reg, col_reg}<13'b1100100110001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b1100100110001) && ({row_reg, col_reg}<13'b1100100110011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1100100110011) && ({row_reg, col_reg}<13'b1100100110111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b1100100110111) && ({row_reg, col_reg}<13'b1100100111001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1100100111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1100100111010) && ({row_reg, col_reg}<13'b1100100111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1100100111110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=13'b1100100111111) && ({row_reg, col_reg}<13'b1100110001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1100110001000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==13'b1100110001001)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==13'b1100110001010)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==13'b1100110001011)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==13'b1100110001100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=13'b1100110001101) && ({row_reg, col_reg}<13'b1100110001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1100110001111) && ({row_reg, col_reg}<13'b1100110010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1100110010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b1100110010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1100110010011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1100110010100) && ({row_reg, col_reg}<13'b1100110010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1100110010111) && ({row_reg, col_reg}<13'b1100110011100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1100110011100) && ({row_reg, col_reg}<13'b1100110100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1100110100110) && ({row_reg, col_reg}<13'b1100110101000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b1100110101000) && ({row_reg, col_reg}<13'b1100110101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1100110101010) && ({row_reg, col_reg}<13'b1100110110111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1100110110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1100110111000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1100110111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1100110111010) && ({row_reg, col_reg}<13'b1100110111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1100110111110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=13'b1100110111111) && ({row_reg, col_reg}<13'b1101000000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1101000000111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==13'b1101000001000)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==13'b1101000001001)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==13'b1101000001010)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==13'b1101000001011)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}>=13'b1101000001100) && ({row_reg, col_reg}<13'b1101000001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b1101000001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1101000001111) && ({row_reg, col_reg}<13'b1101000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1101000010001) && ({row_reg, col_reg}<13'b1101000010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1101000010101) && ({row_reg, col_reg}<13'b1101000011001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1101000011001) && ({row_reg, col_reg}<13'b1101000100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1101000100011) && ({row_reg, col_reg}<13'b1101000101101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1101000101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b1101000101110) && ({row_reg, col_reg}<13'b1101000111001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1101000111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1101000111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1101000111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1101000111100) && ({row_reg, col_reg}<13'b1101000111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1101000111110) && ({row_reg, col_reg}<13'b1101001000000)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=13'b1101001000000) && ({row_reg, col_reg}<13'b1101010000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1101010000110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==13'b1101010000111)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}>=13'b1101010001000) && ({row_reg, col_reg}<13'b1101010001011)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==13'b1101010001011)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}>=13'b1101010001100) && ({row_reg, col_reg}<13'b1101010001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1101010001111) && ({row_reg, col_reg}<13'b1101010010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1101010010101) && ({row_reg, col_reg}<13'b1101010011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1101010011000) && ({row_reg, col_reg}<13'b1101010100010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1101010100010) && ({row_reg, col_reg}<13'b1101010101001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b1101010101001) && ({row_reg, col_reg}<13'b1101010110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b1101010110000) && ({row_reg, col_reg}<13'b1101010111001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1101010111001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1101010111010) && ({row_reg, col_reg}<13'b1101010111101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1101010111101) && ({row_reg, col_reg}<13'b1101010111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1101010111111)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=13'b1101011000000) && ({row_reg, col_reg}<13'b1101100000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1101100000101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b1101100000110)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=13'b1101100000111) && ({row_reg, col_reg}<13'b1101100001011)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==13'b1101100001011)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}>=13'b1101100001100) && ({row_reg, col_reg}<13'b1101100001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1101100001110) && ({row_reg, col_reg}<13'b1101100010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1101100010101) && ({row_reg, col_reg}<13'b1101100010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1101100010111) && ({row_reg, col_reg}<13'b1101100100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1101100100000) && ({row_reg, col_reg}<13'b1101100101000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b1101100101000) && ({row_reg, col_reg}<13'b1101100110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b1101100110000) && ({row_reg, col_reg}<13'b1101100110111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b1101100110111) && ({row_reg, col_reg}<13'b1101100111010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1101100111010) && ({row_reg, col_reg}<13'b1101100111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1101100111111)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=13'b1101101000000) && ({row_reg, col_reg}<13'b1101110000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1101110000100)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==13'b1101110000101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==13'b1101110000110)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==13'b1101110000111)) color_data = 12'b100101100011;
		if(({row_reg, col_reg}==13'b1101110001000)) color_data = 12'b101001100011;
		if(({row_reg, col_reg}==13'b1101110001001)) color_data = 12'b100101100011;
		if(({row_reg, col_reg}==13'b1101110001010)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}>=13'b1101110001011) && ({row_reg, col_reg}<13'b1101110001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1101110001111) && ({row_reg, col_reg}<13'b1101110010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1101110010100) && ({row_reg, col_reg}<13'b1101110011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1101110011000) && ({row_reg, col_reg}<13'b1101110100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1101110100000) && ({row_reg, col_reg}<13'b1101110101000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b1101110101000) && ({row_reg, col_reg}<13'b1101110110001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b1101110110001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b1101110110010) && ({row_reg, col_reg}<13'b1101110110110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b1101110110110) && ({row_reg, col_reg}<13'b1101110111000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1101110111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1101110111001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1101110111010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1101110111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1101110111100) && ({row_reg, col_reg}<13'b1101110111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1101110111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1101110111111) && ({row_reg, col_reg}<13'b1101111000001)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=13'b1101111000001) && ({row_reg, col_reg}<13'b1110000000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1110000000011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b1110000000100)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==13'b1110000000101)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==13'b1110000000110)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==13'b1110000000111)) color_data = 12'b101001100011;
		if(({row_reg, col_reg}==13'b1110000001000)) color_data = 12'b101101110100;
		if(({row_reg, col_reg}==13'b1110000001001)) color_data = 12'b100101100011;
		if(({row_reg, col_reg}==13'b1110000001010)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}>=13'b1110000001011) && ({row_reg, col_reg}<13'b1110000001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1110000001111) && ({row_reg, col_reg}<13'b1110000010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1110000010010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==13'b1110000010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1110000010100) && ({row_reg, col_reg}<13'b1110000011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1110000011000) && ({row_reg, col_reg}<13'b1110000011111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1110000011111) && ({row_reg, col_reg}<13'b1110000100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1110000100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b1110000100100) && ({row_reg, col_reg}<13'b1110000100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b1110000100110) && ({row_reg, col_reg}<13'b1110000110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b1110000110100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1110000110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b1110000110110) && ({row_reg, col_reg}<13'b1110000111000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1110000111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1110000111001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1110000111010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==13'b1110000111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1110000111100) && ({row_reg, col_reg}<13'b1110000111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1110000111110) && ({row_reg, col_reg}<13'b1110001000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1110001000000)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=13'b1110001000001) && ({row_reg, col_reg}<13'b1110010000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1110010000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b1110010000011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==13'b1110010000100)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==13'b1110010000101)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==13'b1110010000110)) color_data = 12'b100101100011;
		if(({row_reg, col_reg}==13'b1110010000111)) color_data = 12'b101101110100;
		if(({row_reg, col_reg}==13'b1110010001000)) color_data = 12'b101001100011;
		if(({row_reg, col_reg}==13'b1110010001001)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==13'b1110010001010)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}>=13'b1110010001011) && ({row_reg, col_reg}<13'b1110010001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1110010001110) && ({row_reg, col_reg}<13'b1110010010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1110010010001) && ({row_reg, col_reg}<13'b1110010011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1110010011000) && ({row_reg, col_reg}<13'b1110010011111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1110010011111) && ({row_reg, col_reg}<13'b1110010100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1110010100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b1110010100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b1110010100101) && ({row_reg, col_reg}<13'b1110010110110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b1110010110110) && ({row_reg, col_reg}<13'b1110010111010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1110010111010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1110010111011) && ({row_reg, col_reg}<13'b1110011000001)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=13'b1110011000001) && ({row_reg, col_reg}<13'b1110100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1110100000001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b1110100000010)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==13'b1110100000011)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==13'b1110100000100)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==13'b1110100000101)) color_data = 12'b101001100011;
		if(({row_reg, col_reg}==13'b1110100000110)) color_data = 12'b101101110100;
		if(({row_reg, col_reg}==13'b1110100000111)) color_data = 12'b110010000101;
		if(({row_reg, col_reg}==13'b1110100001000)) color_data = 12'b101101110100;
		if(({row_reg, col_reg}==13'b1110100001001)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}>=13'b1110100001010) && ({row_reg, col_reg}<13'b1110100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1110100001101) && ({row_reg, col_reg}<13'b1110100001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1110100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b1110100010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1110100010001) && ({row_reg, col_reg}<13'b1110100010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1110100010111) && ({row_reg, col_reg}<13'b1110100011110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1110100011110) && ({row_reg, col_reg}<13'b1110100100010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b1110100100010) && ({row_reg, col_reg}<13'b1110100101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b1110100101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b1110100101111) && ({row_reg, col_reg}<13'b1110100110110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b1110100110110) && ({row_reg, col_reg}<13'b1110100111011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b1110100111011) && ({row_reg, col_reg}<13'b1110101000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1110101000001)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=13'b1110101000010) && ({row_reg, col_reg}<13'b1110110000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1110110000001)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==13'b1110110000010)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==13'b1110110000011)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==13'b1110110000100)) color_data = 12'b101001100011;
		if(({row_reg, col_reg}==13'b1110110000101)) color_data = 12'b101101110100;
		if(({row_reg, col_reg}>=13'b1110110000110) && ({row_reg, col_reg}<13'b1110110001000)) color_data = 12'b110010000101;
		if(({row_reg, col_reg}==13'b1110110001000)) color_data = 12'b101001100011;
		if(({row_reg, col_reg}==13'b1110110001001)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==13'b1110110001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1110110001011) && ({row_reg, col_reg}<13'b1110110001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1110110001101) && ({row_reg, col_reg}<13'b1110110010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1110110010001) && ({row_reg, col_reg}<13'b1110110010110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1110110010110) && ({row_reg, col_reg}<13'b1110110011100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1110110011100) && ({row_reg, col_reg}<13'b1110110100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b1110110100011) && ({row_reg, col_reg}<13'b1110110101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b1110110101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b1110110101100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b1110110101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==13'b1110110101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b1110110101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b1110110110000) && ({row_reg, col_reg}<13'b1110110110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==13'b1110110110101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1110110110110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b1110110110111) && ({row_reg, col_reg}<13'b1110110111011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1110110111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1110110111100) && ({row_reg, col_reg}<13'b1110111000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1110111000001)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}==13'b1110111000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1111000000000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==13'b1111000000001)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}>=13'b1111000000010) && ({row_reg, col_reg}<13'b1111000000100)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==13'b1111000000100)) color_data = 12'b101001100011;
		if(({row_reg, col_reg}==13'b1111000000101)) color_data = 12'b101101110100;
		if(({row_reg, col_reg}==13'b1111000000110)) color_data = 12'b110010000101;
		if(({row_reg, col_reg}==13'b1111000000111)) color_data = 12'b101101110100;
		if(({row_reg, col_reg}==13'b1111000001000)) color_data = 12'b100101100011;
		if(({row_reg, col_reg}==13'b1111000001001)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}>=13'b1111000001010) && ({row_reg, col_reg}<13'b1111000001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1111000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1111000001101) && ({row_reg, col_reg}<13'b1111000010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1111000010001) && ({row_reg, col_reg}<13'b1111000010101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1111000010101) && ({row_reg, col_reg}<13'b1111000011100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1111000011100) && ({row_reg, col_reg}<13'b1111000100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b1111000100100) && ({row_reg, col_reg}<13'b1111000101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b1111000101001) && ({row_reg, col_reg}<13'b1111000110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b1111000110000) && ({row_reg, col_reg}<13'b1111000110111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b1111000110111) && ({row_reg, col_reg}<13'b1111000111011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1111000111011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1111000111100) && ({row_reg, col_reg}<13'b1111001000010)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}==13'b1111001000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==13'b1111010000000)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==13'b1111010000001)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==13'b1111010000010)) color_data = 12'b100101100011;
		if(({row_reg, col_reg}==13'b1111010000011)) color_data = 12'b101001100011;
		if(({row_reg, col_reg}==13'b1111010000100)) color_data = 12'b101101110100;
		if(({row_reg, col_reg}>=13'b1111010000101) && ({row_reg, col_reg}<13'b1111010000111)) color_data = 12'b110010000101;
		if(({row_reg, col_reg}==13'b1111010000111)) color_data = 12'b101001100011;
		if(({row_reg, col_reg}==13'b1111010001000)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}>=13'b1111010001001) && ({row_reg, col_reg}<13'b1111010001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==13'b1111010001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==13'b1111010001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=13'b1111010001101) && ({row_reg, col_reg}<13'b1111010010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=13'b1111010010000) && ({row_reg, col_reg}<13'b1111010010011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=13'b1111010010011) && ({row_reg, col_reg}<13'b1111010011011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1111010011011) && ({row_reg, col_reg}<13'b1111010100001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=13'b1111010100001) && ({row_reg, col_reg}<13'b1111010101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b1111010101011) && ({row_reg, col_reg}<13'b1111010110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=13'b1111010110001) && ({row_reg, col_reg}<13'b1111010111000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=13'b1111010111000) && ({row_reg, col_reg}<13'b1111010111011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==13'b1111010111011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=13'b1111010111100) && ({row_reg, col_reg}<13'b1111011000010)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=13'b1111011000010) && ({row_reg, col_reg}<=13'b1111011000010)) color_data = 12'b000100010001;
	end
endmodule